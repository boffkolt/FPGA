library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use work.lib_lcd.all;
use work.lcd_init.all;

entity LCD is
	
	port( 
		in_std_clk 					:	in std_logic; 	-- тактовая частота	
		in_std_ena					:	in std_logic := '1';														
		out_std7_data				:	out std_logic_vector(7 downto 0) := X"11";
		out_std_cs					:	out std_logic	:= '1';
		out_std_wr					:	out std_logic	:= '1';
		out_std_res					:	out std_logic 	:= '1';
		out_std_a					:	out std_logic 	:= '1';
		out_std_oe_buf				:	out std_logic 	;
		
		out_std_str					:	out std_logic	:= '0';
		in_std_lcd_mode				:	in	std_logic;
		in_std8_data_in				:	in std_logic_vector(7 downto 0) ;
		in_std16_adress				: 	in std_logic_vector(15 downto 0);
		in_std_nwe					:	in	std_logic

	);
		
		
end LCD;
		
architecture LCD_ARCH of LCD is

signal system_set : data (0 to 15) 	:= (	0 	=>	X"40",
															1	=>	X"33",
															2	=>	X"87",
											3	=>	X"07",
											4	=>	X"27",
											5	=>	X"2F",
											6	=>	X"EF",
											7	=>	X"28",
											8	=>	X"00",
											others=> X"00");
								
								
signal scroll : data (0 to 15)		:= (0	=>	X"44",
											1	=>	X"00",
											2	=>	X"00",
											3	=>	X"EF",
											4	=>	X"B0",
											5	=>	X"04",
											6	=>	X"EF",
											7	=>	X"30",
											8	=>	X"2A",
											9	=>	X"00",
											10	=>	X"00",
											others=> X"00");
								
signal hdot_scr : data (0 to 1)		:= (0	=>	X"5A",
												1	=>	X"00");
								
signal ovlay : data (0 to 1)			:= (0	=>	X"5B",
											1	=>	X"01");

signal cgram_adr : data (0 to 3)		:= (0	=>	X"5C",
											1	=>	X"00",
											2	=> X"F0",
											others=> X"00");
											
signal disp_off : data (0 to 1)		:= (0	=>	X"58",
											1	=>	X"56");
											
signal disp_on : data (0 to 1)		:= (0	=>	X"59",
											1	=>	X"10");
											
signal set_start_clr : data (0 to 3)	:= (0	=>	X"46",
											1	=>	X"00",
											2 	=>	X"00",
											others=> X"00");
											
signal set_start : data (0 to 3)		:= (0	=>	X"46",
											1	=>	X"B0",
											2 	=>	X"04",
											others=> X"00");
											
signal clr_disp : data (0 to 16383)	:= (	0	=>	X"42",
											others	=>	X"00");	
											
signal logo_elsiel : data (0 to 16383) 	:= (	0 	=> X"42",
																1	=> X"00",
																2	=>	X"00",
																3	=>	X"00",
																4	=>	X"00",
																5	=>	X"00",
																6	=>	X"00",
																7	=>	X"00",
																8	=>	X"00",
																9	=>	X"00",
																10	=>	X"00",
																11	=>	X"00",
																12	=>	X"00",
																13	=>	X"00",
																14	=>	X"00",
																15	=>	X"00",
																16	=>	X"00",
																17	=>	X"00",
																18	=>	X"00",
																19	=>	X"00",
																20	=>	X"00",
																21	=>	X"00",
																22	=>	X"00",
																23	=>	X"00",
																24	=>	X"00",
																25	=>	X"00",
																26	=>	X"00",
																27	=>	X"00",
																28	=>	X"00",
																29	=>	X"00",
																30	=>	X"00",
																31	=>	X"00",
																32	=>	X"00",
																33	=>	X"00",
																34	=>	X"00",
																35	=>	X"00",
																36	=>	X"00",
																37	=>	X"00",
																38	=>	X"00",
																39	=>	X"00",
																40	=>	X"00",
																41	=>	X"00",
																42	=>	X"00",
																43	=>	X"00",
																44	=>	X"00",
																45	=>	X"00",
																46	=>	X"00",
																47	=>	X"00",
																48	=>	X"00",
																49	=>	X"00",
																50	=>	X"00",
																51	=>	X"00",
																52	=>	X"00",
																53	=>	X"00",
																54	=>	X"00",
																55	=>	X"00",
																56	=>	X"00",
																57	=>	X"00",
																58	=>	X"00",
																59	=>	X"00",
																60	=>	X"00",
																61	=>	X"00",
																62	=>	X"00",
																63	=>	X"00",
																64	=>	X"00",
																65	=>	X"00",
																66	=>	X"00",
																67	=>	X"00",
																68	=>	X"00",
																69	=>	X"00",
																70	=>	X"00",
																71	=>	X"00",
																72	=>	X"00",
																73	=>	X"00",
																74	=>	X"00",
																75	=>	X"00",
																76	=>	X"00",
																77	=>	X"00",
																78	=>	X"00",
																79	=>	X"00",
																80	=>	X"00",
																81	=>	X"00",
																82	=>	X"00",
																83	=>	X"00",
																84	=>	X"00",
																85	=>	X"00",
																86	=>	X"00",
																87	=>	X"00",
																88	=>	X"00",
																89	=>	X"00",
																90	=>	X"00",
																91	=>	X"00",
																92	=>	X"00",
																93	=>	X"00",
																94	=>	X"00",
																95	=>	X"00",
																96	=>	X"00",
																97	=>	X"00",
																98	=>	X"00",
																99	=>	X"00",
																100	=>	X"00",
																101	=>	X"00",
																102	=>	X"00",
																103	=>	X"00",
																104	=>	X"00",
																105	=>	X"00",
																106	=>	X"00",
																107	=>	X"00",
																108	=>	X"00",
																109	=>	X"00",
																110	=>	X"00",
																111	=>	X"00",
																112	=>	X"00",
																113	=>	X"00",
																114	=>	X"00",
																115	=>	X"00",
																116	=>	X"00",
																117	=>	X"00",
																118	=>	X"00",
																119	=>	X"00",
																120	=>	X"00",
																121	=>	X"00",
																122	=>	X"00",
																123	=>	X"00",
																124	=>	X"00",
																125	=>	X"00",
																126	=>	X"00",
																127	=>	X"00",
																128	=>	X"00",
																129	=>	X"00",
																130	=>	X"00",
																131	=>	X"00",
																132	=>	X"00",
																133	=>	X"00",
																134	=>	X"00",
																135	=>	X"00",
																136	=>	X"00",
																137	=>	X"00",
																138	=>	X"00",
																139	=>	X"00",
																140	=>	X"00",
																141	=>	X"00",
																142	=>	X"00",
																143	=>	X"00",
																144	=>	X"00",
																145	=>	X"00",
																146	=>	X"00",
																147	=>	X"00",
																148	=>	X"00",
																149	=>	X"00",
																150	=>	X"00",
																151	=>	X"00",
																152	=>	X"00",
																153	=>	X"00",
																154	=>	X"00",
																155	=>	X"00",
																156	=>	X"00",
																157	=>	X"00",
																158	=>	X"00",
																159	=>	X"00",
																160	=>	X"00",
																161	=>	X"00",
																162	=>	X"00",
																163	=>	X"00",
																164	=>	X"00",
																165	=>	X"00",
																166	=>	X"00",
																167	=>	X"00",
																168	=>	X"00",
																169	=>	X"00",
																170	=>	X"00",
																171	=>	X"00",
																172	=>	X"00",
																173	=>	X"00",
																174	=>	X"00",
																175	=>	X"00",
																176	=>	X"00",
																177	=>	X"00",
																178	=>	X"00",
																179	=>	X"00",
																180	=>	X"00",
																181	=>	X"00",
																182	=>	X"00",
																183	=>	X"00",
																184	=>	X"00",
																185	=>	X"00",
																186	=>	X"00",
																187	=>	X"00",
																188	=>	X"00",
																189	=>	X"00",
																190	=>	X"00",
																191	=>	X"00",
																192	=>	X"00",
																193	=>	X"00",
																194	=>	X"00",
																195	=>	X"00",
																196	=>	X"00",
																197	=>	X"00",
																198	=>	X"00",
																199	=>	X"00",
																200	=>	X"00",
																201	=>	X"00",
																202	=>	X"00",
																203	=>	X"00",
																204	=>	X"00",
																205	=>	X"00",
																206	=>	X"00",
																207	=>	X"00",
																208	=>	X"00",
																209	=>	X"00",
																210	=>	X"00",
																211	=>	X"00",
																212	=>	X"00",
																213	=>	X"00",
																214	=>	X"00",
																215	=>	X"00",
																216	=>	X"00",
																217	=>	X"00",
																218	=>	X"00",
																219	=>	X"00",
																220	=>	X"00",
																221	=>	X"00",
																222	=>	X"00",
																223	=>	X"00",
																224	=>	X"00",
																225	=>	X"00",
																226	=>	X"00",
																227	=>	X"00",
																228	=>	X"00",
																229	=>	X"00",
																230	=>	X"00",
																231	=>	X"00",
																232	=>	X"00",
																233	=>	X"00",
																234	=>	X"00",
																235	=>	X"00",
																236	=>	X"00",
																237	=>	X"00",
																238	=>	X"00",
																239	=>	X"00",
																240	=>	X"00",
																241	=>	X"00",
																242	=>	X"00",
																243	=>	X"00",
																244	=>	X"00",
																245	=>	X"00",
																246	=>	X"00",
																247	=>	X"00",
																248	=>	X"00",
																249	=>	X"00",
																250	=>	X"00",
																251	=>	X"00",
																252	=>	X"00",
																253	=>	X"00",
																254	=>	X"00",
																255	=>	X"00",
																256	=>	X"00",
																257	=>	X"00",
																258	=>	X"00",
																259	=>	X"00",
																260	=>	X"00",
																261	=>	X"00",
																262	=>	X"00",
																263	=>	X"00",
																264	=>	X"00",
																265	=>	X"00",
																266	=>	X"00",
																267	=>	X"00",
																268	=>	X"00",
																269	=>	X"00",
																270	=>	X"00",
																271	=>	X"00",
																272	=>	X"00",
																273	=>	X"00",
																274	=>	X"00",
																275	=>	X"00",
																276	=>	X"00",
																277	=>	X"00",
																278	=>	X"00",
																279	=>	X"00",
																280	=>	X"00",
																281	=>	X"00",
																282	=>	X"00",
																283	=>	X"00",
																284	=>	X"00",
																285	=>	X"00",
																286	=>	X"00",
																287	=>	X"00",
																288	=>	X"00",
																289	=>	X"00",
																290	=>	X"00",
																291	=>	X"00",
																292	=>	X"00",
																293	=>	X"00",
																294	=>	X"00",
																295	=>	X"00",
																296	=>	X"00",
																297	=>	X"00",
																298	=>	X"00",
																299	=>	X"00",
																300	=>	X"00",
																301	=>	X"00",
																302	=>	X"00",
																303	=>	X"00",
																304	=>	X"00",
																305	=>	X"00",
																306	=>	X"00",
																307	=>	X"00",
																308	=>	X"00",
																309	=>	X"00",
																310	=>	X"00",
																311	=>	X"00",
																312	=>	X"00",
																313	=>	X"00",
																314	=>	X"00",
																315	=>	X"00",
																316	=>	X"00",
																317	=>	X"00",
																318	=>	X"00",
																319	=>	X"00",
																320	=>	X"00",
																321	=>	X"00",
																322	=>	X"00",
																323	=>	X"00",
																324	=>	X"00",
																325	=>	X"00",
																326	=>	X"00",
																327	=>	X"00",
																328	=>	X"00",
																329	=>	X"00",
																330	=>	X"00",
																331	=>	X"00",
																332	=>	X"00",
																333	=>	X"00",
																334	=>	X"00",
																335	=>	X"00",
																336	=>	X"00",
																337	=>	X"00",
																338	=>	X"00",
																339	=>	X"00",
																340	=>	X"00",
																341	=>	X"00",
																342	=>	X"00",
																343	=>	X"00",
																344	=>	X"00",
																345	=>	X"00",
																346	=>	X"00",
																347	=>	X"00",
																348	=>	X"00",
																349	=>	X"00",
																350	=>	X"00",
																351	=>	X"00",
																352	=>	X"00",
																353	=>	X"00",
																354	=>	X"00",
																355	=>	X"00",
																356	=>	X"00",
																357	=>	X"00",
																358	=>	X"00",
																359	=>	X"00",
																360	=>	X"00",
																361	=>	X"00",
																362	=>	X"00",
																363	=>	X"00",
																364	=>	X"00",
																365	=>	X"00",
																366	=>	X"00",
																367	=>	X"00",
																368	=>	X"00",
																369	=>	X"00",
																370	=>	X"00",
																371	=>	X"00",
																372	=>	X"00",
																373	=>	X"00",
																374	=>	X"00",
																375	=>	X"00",
																376	=>	X"00",
																377	=>	X"00",
																378	=>	X"00",
																379	=>	X"00",
																380	=>	X"00",
																381	=>	X"00",
																382	=>	X"00",
																383	=>	X"00",
																384	=>	X"00",
																385	=>	X"00",
																386	=>	X"00",
																387	=>	X"00",
																388	=>	X"00",
																389	=>	X"00",
																390	=>	X"00",
																391	=>	X"00",
																392	=>	X"00",
																393	=>	X"00",
																394	=>	X"00",
																395	=>	X"00",
																396	=>	X"00",
																397	=>	X"00",
																398	=>	X"00",
																399	=>	X"00",
																400	=>	X"00",
																401	=>	X"00",
																402	=>	X"00",
																403	=>	X"00",
																404	=>	X"00",
																405	=>	X"00",
																406	=>	X"00",
																407	=>	X"00",
																408	=>	X"00",
																409	=>	X"00",
																410	=>	X"00",
																411	=>	X"00",
																412	=>	X"00",
																413	=>	X"00",
																414	=>	X"00",
																415	=>	X"00",
																416	=>	X"00",
																417	=>	X"00",
																418	=>	X"00",
																419	=>	X"00",
																420	=>	X"00",
																421	=>	X"00",
																422	=>	X"00",
																423	=>	X"00",
																424	=>	X"00",
																425	=>	X"00",
																426	=>	X"00",
																427	=>	X"00",
																428	=>	X"00",
																429	=>	X"00",
																430	=>	X"00",
																431	=>	X"00",
																432	=>	X"00",
																433	=>	X"00",
																434	=>	X"00",
																435	=>	X"00",
																436	=>	X"00",
																437	=>	X"00",
																438	=>	X"00",
																439	=>	X"00",
																440	=>	X"00",
																441	=>	X"00",
																442	=>	X"00",
																443	=>	X"00",
																444	=>	X"00",
																445	=>	X"00",
																446	=>	X"00",
																447	=>	X"00",
																448	=>	X"00",
																449	=>	X"00",
																450	=>	X"00",
																451	=>	X"00",
																452	=>	X"00",
																453	=>	X"00",
																454	=>	X"00",
																455	=>	X"00",
																456	=>	X"00",
																457	=>	X"00",
																458	=>	X"00",
																459	=>	X"00",
																460	=>	X"00",
																461	=>	X"00",
																462	=>	X"00",
																463	=>	X"00",
																464	=>	X"00",
																465	=>	X"00",
																466	=>	X"00",
																467	=>	X"00",
																468	=>	X"00",
																469	=>	X"00",
																470	=>	X"00",
																471	=>	X"00",
																472	=>	X"00",
																473	=>	X"00",
																474	=>	X"00",
																475	=>	X"00",
																476	=>	X"00",
																477	=>	X"00",
																478	=>	X"00",
																479	=>	X"00",
																480	=>	X"00",
																481	=>	X"00",
																482	=>	X"00",
																483	=>	X"00",
																484	=>	X"00",
																485	=>	X"00",
																486	=>	X"00",
																487	=>	X"00",
																488	=>	X"00",
																489	=>	X"00",
																490	=>	X"00",
																491	=>	X"00",
																492	=>	X"00",
																493	=>	X"00",
																494	=>	X"00",
																495	=>	X"00",
																496	=>	X"00",
																497	=>	X"00",
																498	=>	X"00",
																499	=>	X"00",
																500	=>	X"00",
																501	=>	X"00",
																502	=>	X"00",
																503	=>	X"00",
																504	=>	X"00",
																505	=>	X"00",
																506	=>	X"00",
																507	=>	X"00",
																508	=>	X"00",
																509	=>	X"00",
																510	=>	X"00",
																511	=>	X"00",
																512	=>	X"00",
																513	=>	X"00",
																514	=>	X"00",
																515	=>	X"00",
																516	=>	X"00",
																517	=>	X"00",
																518	=>	X"00",
																519	=>	X"00",
																520	=>	X"00",
																521	=>	X"00",
																522	=>	X"00",
																523	=>	X"00",
																524	=>	X"00",
																525	=>	X"00",
																526	=>	X"00",
																527	=>	X"00",
																528	=>	X"00",
																529	=>	X"00",
																530	=>	X"00",
																531	=>	X"00",
																532	=>	X"00",
																533	=>	X"00",
																534	=>	X"00",
																535	=>	X"00",
																536	=>	X"00",
																537	=>	X"00",
																538	=>	X"00",
																539	=>	X"00",
																540	=>	X"00",
																541	=>	X"00",
																542	=>	X"00",
																543	=>	X"00",
																544	=>	X"00",
																545	=>	X"00",
																546	=>	X"00",
																547	=>	X"00",
																548	=>	X"00",
																549	=>	X"00",
																550	=>	X"00",
																551	=>	X"00",
																552	=>	X"00",
																553	=>	X"00",
																554	=>	X"00",
																555	=>	X"00",
																556	=>	X"00",
																557	=>	X"00",
																558	=>	X"00",
																559	=>	X"00",
																560	=>	X"00",
																561	=>	X"00",
																562	=>	X"00",
																563	=>	X"00",
																564	=>	X"00",
																565	=>	X"00",
																566	=>	X"00",
																567	=>	X"00",
																568	=>	X"00",
																569	=>	X"00",
																570	=>	X"00",
																571	=>	X"00",
																572	=>	X"00",
																573	=>	X"00",
																574	=>	X"00",
																575	=>	X"00",
																576	=>	X"00",
																577	=>	X"00",
																578	=>	X"00",
																579	=>	X"00",
																580	=>	X"00",
																581	=>	X"00",
																582	=>	X"00",
																583	=>	X"00",
																584	=>	X"00",
																585	=>	X"00",
																586	=>	X"00",
																587	=>	X"00",
																588	=>	X"00",
																589	=>	X"00",
																590	=>	X"00",
																591	=>	X"00",
																592	=>	X"00",
																593	=>	X"00",
																594	=>	X"00",
																595	=>	X"00",
																596	=>	X"00",
																597	=>	X"00",
																598	=>	X"00",
																599	=>	X"00",
																600	=>	X"00",
																601	=>	X"00",
																602	=>	X"00",
																603	=>	X"00",
																604	=>	X"00",
																605	=>	X"00",
																606	=>	X"00",
																607	=>	X"00",
																608	=>	X"00",
																609	=>	X"00",
																610	=>	X"00",
																611	=>	X"00",
																612	=>	X"00",
																613	=>	X"00",
																614	=>	X"00",
																615	=>	X"00",
																616	=>	X"00",
																617	=>	X"00",
																618	=>	X"00",
																619	=>	X"00",
																620	=>	X"00",
																621	=>	X"00",
																622	=>	X"00",
																623	=>	X"00",
																624	=>	X"00",
																625	=>	X"00",
																626	=>	X"00",
																627	=>	X"00",
																628	=>	X"00",
																629	=>	X"00",
																630	=>	X"00",
																631	=>	X"00",
																632	=>	X"00",
																633	=>	X"00",
																634	=>	X"00",
																635	=>	X"00",
																636	=>	X"00",
																637	=>	X"00",
																638	=>	X"00",
																639	=>	X"00",
																640	=>	X"00",
																641	=>	X"00",
																642	=>	X"00",
																643	=>	X"00",
																644	=>	X"00",
																645	=>	X"00",
																646	=>	X"00",
																647	=>	X"00",
																648	=>	X"00",
																649	=>	X"00",
																650	=>	X"00",
																651	=>	X"00",
																652	=>	X"00",
																653	=>	X"00",
																654	=>	X"00",
																655	=>	X"00",
																656	=>	X"00",
																657	=>	X"00",
																658	=>	X"00",
																659	=>	X"00",
																660	=>	X"00",
																661	=>	X"00",
																662	=>	X"00",
																663	=>	X"00",
																664	=>	X"00",
																665	=>	X"00",
																666	=>	X"00",
																667	=>	X"00",
																668	=>	X"00",
																669	=>	X"00",
																670	=>	X"00",
																671	=>	X"00",
																672	=>	X"00",
																673	=>	X"00",
																674	=>	X"00",
																675	=>	X"00",
																676	=>	X"00",
																677	=>	X"00",
																678	=>	X"00",
																679	=>	X"00",
																680	=>	X"00",
																681	=>	X"00",
																682	=>	X"00",
																683	=>	X"00",
																684	=>	X"00",
																685	=>	X"00",
																686	=>	X"00",
																687	=>	X"00",
																688	=>	X"00",
																689	=>	X"00",
																690	=>	X"00",
																691	=>	X"00",
																692	=>	X"00",
																693	=>	X"00",
																694	=>	X"00",
																695	=>	X"00",
																696	=>	X"00",
																697	=>	X"00",
																698	=>	X"00",
																699	=>	X"00",
																700	=>	X"00",
																701	=>	X"00",
																702	=>	X"00",
																703	=>	X"00",
																704	=>	X"00",
																705	=>	X"00",
																706	=>	X"00",
																707	=>	X"00",
																708	=>	X"00",
																709	=>	X"00",
																710	=>	X"00",
																711	=>	X"00",
																712	=>	X"00",
																713	=>	X"00",
																714	=>	X"00",
																715	=>	X"00",
																716	=>	X"00",
																717	=>	X"00",
																718	=>	X"00",
																719	=>	X"00",
																720	=>	X"00",
																721	=>	X"00",
																722	=>	X"00",
																723	=>	X"00",
																724	=>	X"00",
																725	=>	X"00",
																726	=>	X"00",
																727	=>	X"00",
																728	=>	X"00",
																729	=>	X"00",
																730	=>	X"00",
																731	=>	X"00",
																732	=>	X"00",
																733	=>	X"00",
																734	=>	X"00",
																735	=>	X"00",
																736	=>	X"00",
																737	=>	X"00",
																738	=>	X"00",
																739	=>	X"00",
																740	=>	X"00",
																741	=>	X"00",
																742	=>	X"00",
																743	=>	X"00",
																744	=>	X"00",
																745	=>	X"00",
																746	=>	X"00",
																747	=>	X"00",
																748	=>	X"00",
																749	=>	X"00",
																750	=>	X"00",
																751	=>	X"00",
																752	=>	X"00",
																753	=>	X"00",
																754	=>	X"00",
																755	=>	X"00",
																756	=>	X"00",
																757	=>	X"00",
																758	=>	X"00",
																759	=>	X"00",
																760	=>	X"00",
																761	=>	X"00",
																762	=>	X"00",
																763	=>	X"00",
																764	=>	X"00",
																765	=>	X"00",
																766	=>	X"00",
																767	=>	X"00",
																768	=>	X"00",
																769	=>	X"00",
																770	=>	X"00",
																771	=>	X"00",
																772	=>	X"00",
																773	=>	X"00",
																774	=>	X"00",
																775	=>	X"00",
														776	=>	X"00",
														777	=>	X"00",
														778	=>	X"00",
														779	=>	X"00",
														780	=>	X"00",
														781	=>	X"00",
														782	=>	X"00",
														783	=>	X"00",
														784	=>	X"00",
														785	=>	X"00",
														786	=>	X"00",
														787	=>	X"00",
														788	=>	X"00",
														789	=>	X"00",
														790	=>	X"00",
														791	=>	X"00",
														792	=>	X"00",
														793	=>	X"00",
														794	=>	X"00",
														795	=>	X"00",
														796	=>	X"00",
														797	=>	X"00",
														798	=>	X"00",
														799	=>	X"00",
														800	=>	X"00",
														801	=>	X"00",
														802	=>	X"00",
														803	=>	X"00",
														804	=>	X"00",
														805	=>	X"00",
														806	=>	X"00",
														807	=>	X"00",
														808	=>	X"00",
														809	=>	X"00",
														810	=>	X"00",
														811	=>	X"00",
														812	=>	X"00",
														813	=>	X"00",
														814	=>	X"00",
														815	=>	X"00",
														816	=>	X"00",
														817	=>	X"00",
														818	=>	X"00",
														819	=>	X"00",
														820	=>	X"00",
														821	=>	X"00",
														822	=>	X"00",
														823	=>	X"00",
														824	=>	X"00",
														825	=>	X"00",
														826	=>	X"00",
														827	=>	X"00",
														828	=>	X"00",
														829	=>	X"00",
														830	=>	X"00",
														831	=>	X"00",
														832	=>	X"00",
														833	=>	X"00",
														834	=>	X"00",
														835	=>	X"00",
														836	=>	X"00",
														837	=>	X"00",
														838	=>	X"00",
														839	=>	X"00",
														840	=>	X"00",
														841	=>	X"00",
														842	=>	X"00",
														843	=>	X"00",
														844	=>	X"00",
														845	=>	X"00",
														846	=>	X"00",
														847	=>	X"00",
														848	=>	X"00",
														849	=>	X"00",
														850	=>	X"00",
														851	=>	X"00",
														852	=>	X"00",
														853	=>	X"00",
														854	=>	X"00",
														855	=>	X"00",
														856	=>	X"00",
														857	=>	X"00",
														858	=>	X"00",
														859	=>	X"00",
														860	=>	X"00",
														861	=>	X"00",
														862	=>	X"00",
														863	=>	X"00",
														864	=>	X"00",
														865	=>	X"00",
														866	=>	X"00",
														867	=>	X"00",
														868	=>	X"00",
														869	=>	X"00",
														870	=>	X"00",
														871	=>	X"00",
														872	=>	X"00",
														873	=>	X"00",
														874	=>	X"00",
														875	=>	X"00",
														876	=>	X"00",
														877	=>	X"00",
														878	=>	X"00",
														879	=>	X"00",
														880	=>	X"00",
														881	=>	X"00",
														882	=>	X"00",
														883	=>	X"00",
														884	=>	X"00",
														885	=>	X"00",
														886	=>	X"00",
														887	=>	X"00",
														888	=>	X"00",
														889	=>	X"00",
														890	=>	X"00",
														891	=>	X"00",
														892	=>	X"00",
														893	=>	X"00",
														894	=>	X"00",
														895	=>	X"00",
														896	=>	X"00",
														897	=>	X"00",
														898	=>	X"00",
														899	=>	X"00",
														900	=>	X"00",
														901	=>	X"00",
														902	=>	X"00",
														903	=>	X"00",
														904	=>	X"00",
														905	=>	X"00",
														906	=>	X"00",
														907	=>	X"00",
														908	=>	X"00",
														909	=>	X"00",
														910	=>	X"00",
														911	=>	X"00",
														912	=>	X"00",
														913	=>	X"00",
														914	=>	X"00",
														915	=>	X"00",
														916	=>	X"00",
														917	=>	X"00",
														918	=>	X"00",
														919	=>	X"00",
														920	=>	X"00",
														921	=>	X"00",
														922	=>	X"00",
														923	=>	X"00",
														924	=>	X"00",
														925	=>	X"00",
														926	=>	X"00",
														927	=>	X"00",
														928	=>	X"00",
														929	=>	X"00",
														930	=>	X"00",
														931	=>	X"00",
														932	=>	X"00",
														933	=>	X"00",
														934	=>	X"00",
														935	=>	X"00",
														936	=>	X"00",
														937	=>	X"00",
														938	=>	X"00",
														939	=>	X"00",
														940	=>	X"00",
														941	=>	X"00",
														942	=>	X"00",
														943	=>	X"00",
														944	=>	X"00",
														945	=>	X"00",
														946	=>	X"00",
														947	=>	X"00",
														948	=>	X"00",
														949	=>	X"00",
														950	=>	X"00",
														951	=>	X"00",
														952	=>	X"00",
														953	=>	X"00",
														954	=>	X"00",
														955	=>	X"00",
														956	=>	X"00",
														957	=>	X"00",
														958	=>	X"00",
														959	=>	X"00",
														960	=>	X"00",
														961	=>	X"00",
														962	=>	X"00",
														963	=>	X"00",
														964	=>	X"00",
														965	=>	X"00",
														966	=>	X"00",
														967	=>	X"00",
														968	=>	X"00",
														969	=>	X"00",
														970	=>	X"00",
														971	=>	X"00",
														972	=>	X"00",
														973	=>	X"00",
														974	=>	X"00",
														975	=>	X"00",
														976	=>	X"00",
														977	=>	X"00",
														978	=>	X"00",
														979	=>	X"00",
														980	=>	X"00",
														981	=>	X"00",
														982	=>	X"00",
														983	=>	X"00",
														984	=>	X"00",
														985	=>	X"00",
														986	=>	X"00",
														987	=>	X"00",
														988	=>	X"00",
														989	=>	X"00",
														990	=>	X"00",
														991	=>	X"00",
														992	=>	X"00",
														993	=>	X"00",
														994	=>	X"00",
														995	=>	X"00",
														996	=>	X"00",
														997	=>	X"00",
														998	=>	X"00",
														999	=>	X"00",
														1000	=>	X"00",
														1001	=>	X"00",
														1002	=>	X"00",
														1003	=>	X"00",
														1004	=>	X"00",
														1005	=>	X"00",
														1006	=>	X"00",
														1007	=>	X"00",
														1008	=>	X"00",
														1009	=>	X"00",
														1010	=>	X"00",
														1011	=>	X"00",
														1012	=>	X"00",
														1013	=>	X"00",
														1014	=>	X"00",
														1015	=>	X"00",
														1016	=>	X"00",
														1017	=>	X"00",
														1018	=>	X"00",
														1019	=>	X"00",
														1020	=>	X"00",
														1021	=>	X"00",
														1022	=>	X"00",
														1023	=>	X"00",
														1024	=>	X"00",
														1025	=>	X"00",
														1026	=>	X"00",
														1027	=>	X"00",
														1028	=>	X"00",
														1029	=>	X"00",
														1030	=>	X"00",
														1031	=>	X"00",
														1032	=>	X"00",
														1033	=>	X"00",
														1034	=>	X"00",
														1035	=>	X"00",
														1036	=>	X"00",
														1037	=>	X"00",
														1038	=>	X"00",
														1039	=>	X"00",
														1040	=>	X"00",
														1041	=>	X"00",
														1042	=>	X"00",
														1043	=>	X"00",
														1044	=>	X"00",
														1045	=>	X"00",
														1046	=>	X"00",
														1047	=>	X"00",
														1048	=>	X"00",
														1049	=>	X"00",
														1050	=>	X"00",
														1051	=>	X"00",
														1052	=>	X"00",
														1053	=>	X"00",
														1054	=>	X"00",
														1055	=>	X"00",
														1056	=>	X"00",
														1057	=>	X"00",
														1058	=>	X"00",
														1059	=>	X"00",
														1060	=>	X"00",
														1061	=>	X"00",
														1062	=>	X"00",
														1063	=>	X"00",
														1064	=>	X"00",
														1065	=>	X"00",
														1066	=>	X"00",
														1067	=>	X"00",
														1068	=>	X"00",
														1069	=>	X"00",
														1070	=>	X"00",
														1071	=>	X"00",
														1072	=>	X"00",
														1073	=>	X"00",
														1074	=>	X"00",
														1075	=>	X"00",
														1076	=>	X"00",
														1077	=>	X"00",
														1078	=>	X"00",
														1079	=>	X"00",
														1080	=>	X"00",
														1081	=>	X"00",
														1082	=>	X"00",
														1083	=>	X"00",
														1084	=>	X"00",
														1085	=>	X"00",
														1086	=>	X"00",
														1087	=>	X"00",
														1088	=>	X"00",
														1089	=>	X"00",
														1090	=>	X"00",
														1091	=>	X"00",
														1092	=>	X"00",
														1093	=>	X"00",
														1094	=>	X"00",
														1095	=>	X"00",
														1096	=>	X"00",
														1097	=>	X"00",
														1098	=>	X"00",
														1099	=>	X"00",
														1100	=>	X"00",
														1101	=>	X"00",
														1102	=>	X"00",
														1103	=>	X"00",
														1104	=>	X"00",
														1105	=>	X"00",
														1106	=>	X"00",
														1107	=>	X"00",
														1108	=>	X"00",
														1109	=>	X"00",
														1110	=>	X"00",
														1111	=>	X"00",
														1112	=>	X"00",
														1113	=>	X"00",
														1114	=>	X"00",
														1115	=>	X"00",
														1116	=>	X"00",
														1117	=>	X"00",
														1118	=>	X"00",
														1119	=>	X"00",
														1120	=>	X"00",
														1121	=>	X"00",
														1122	=>	X"00",
														1123	=>	X"00",
														1124	=>	X"00",
														1125	=>	X"00",
														1126	=>	X"00",
														1127	=>	X"00",
													1128	=>X"00",
													1129	=>X"00",
													1130	=>X"00",
													1131	=>X"00",
													1132	=>X"00",
													1133	=>X"00",
													1134	=>X"00",
													1135	=>X"00",
													1136	=>X"00",
													1137	=>X"00",
													1138	=>X"00",
													1139	=>X"00",
													1140	=>X"00",
													1141	=>X"00",
													1142	=>X"00",
													1143	=>X"00",
													1144	=>X"00",
													1145	=>X"00",
													1146	=>X"00",
													1147	=>X"00",
													1148	=>X"00",
													1149	=>X"00",
													1150	=>X"00",
													1151	=>X"00",
													1152	=>X"00",
													1153	=>X"00",
													1154	=>X"00",
													1155	=>X"00",
													1156	=>X"00",
													1157	=>X"00",
													1158	=>X"00",
													1159	=>X"00",
													1160	=>X"00",
													1161	=>X"00",
													1162	=>X"00",
													1163	=>X"00",
													1164	=>X"00",
													1165	=>X"00",
													1166	=>X"00",
													1167	=>X"00",
													1168	=>X"00",
													1169	=>X"00",
													1170	=>X"00",
													1171	=>X"00",
													1172	=>X"00",
													1173	=>X"00",
													1174	=>X"00",
													1175	=>X"00",
													1176	=>X"00",
													1177	=>X"00",
													1178	=>X"00",
													1179	=>X"00",
													1180	=>X"00",
													1181	=>X"00",
													1182	=>X"00",
													1183	=>X"00",
													1184	=>X"00",
													1185	=>X"00",
													1186	=>X"00",
													1187	=>X"00",
													1188	=>X"00",
													1189	=>X"00",
													1190	=>X"00",
													1191	=>X"00",
													1192	=>X"00",
													1193	=>X"00",
													1194	=>X"00",
													1195	=>X"00",
													1196	=>X"00",
													1197	=>X"00",
													1198	=>X"00",
													1199	=>X"00",
													1200	=>X"00",
													1201	=>X"00",
													1202	=>X"00",
													1203	=>X"00",
													1204	=>X"00",
													1205	=>X"00",
													1206	=>X"00",
													1207	=>X"00",
													1208	=>X"00",
													1209	=>X"00",
													1210	=>X"00",
													1211	=>X"00",
													1212	=>X"00",
													1213	=>X"00",
													1214	=>X"00",
													1215	=>X"00",
													1216	=>X"00",
													1217	=>X"00",
													1218	=>X"00",
													1219	=>X"00",
													1220	=>X"00",
													1221	=>X"00",
													1222	=>X"00",
													1223	=>X"00",
													1224	=>X"00",
													1225	=>X"00",
													1226	=>X"00",
													1227	=>X"00",
													1228	=>X"00",
													1229	=>X"00",
													1230	=>X"00",
													1231	=>X"00",
													1232	=>X"00",
													1233	=>X"00",
													1234	=>X"00",
													1235	=>X"00",
													1236	=>X"00",
													1237	=>X"00",
													1238	=>X"00",
													1239	=>X"00",
													1240	=>X"00",
													1241	=>X"00",
													1242	=>X"00",
													1243	=>X"00",
													1244	=>X"00",
													1245	=>X"00",
													1246	=>X"00",
													1247	=>X"00",
													1248	=>X"00",
													1249	=>X"00",
													1250	=>X"00",
													1251	=>X"00",
													1252	=>X"00",
													1253	=>X"00",
													1254	=>X"00",
													1255	=>X"00",
													1256	=>X"00",
													1257	=>X"00",
													1258	=>X"00",
													1259	=>X"00",
													1260	=>X"00",
													1261	=>X"00",
													1262	=>X"00",
													1263	=>X"00",
													1264	=>X"00",
													1265	=>X"00",
													1266	=>X"00",
													1267	=>X"00",
													1268	=>X"00",
													1269	=>X"00",
													1270	=>X"00",
													1271	=>X"00",
													1272	=>X"00",
													1273	=>X"00",
													1274	=>X"00",
													1275	=>X"00",
													1276	=>X"00",
													1277	=>X"00",
													1278	=>X"00",
													1279	=>X"00",
													1280	=>X"00",
													1281	=>X"00",
													1282	=>X"00",
													1283	=>X"00",
													1284	=>X"00",
													1285	=>X"00",
													1286	=>X"00",
													1287	=>X"00",
													1288	=>X"00",
													1289	=>X"00",
													1290	=>X"00",
													1291	=>X"00",
													1292	=>X"00",
													1293	=>X"00",
													1294	=>X"00",
													1295	=>X"00",
													1296	=>X"00",
													1297	=>X"00",
													1298	=>X"00",
													1299	=>X"00",
													1300	=>X"00",
													1301	=>X"00",
													1302	=>X"00",
													1303	=>X"00",
													1304	=>X"00",
													1305	=>X"00",
													1306	=>X"00",
													1307	=>X"00",
													1308	=>X"00",
													1309	=>X"00",
													1310	=>X"00",
													1311	=>X"00",
													1312	=>X"00",
													1313	=>X"00",
													1314	=>X"00",
													1315	=>X"00",
													1316	=>X"00",
													1317	=>X"00",
													1318	=>X"00",
													1319	=>X"00",
													1320	=>X"00",
													1321	=>X"00",
													1322	=>X"00",
													1323	=>X"00",
													1324	=>X"00",
													1325	=>X"00",
													1326	=>X"00",
													1327	=>X"00",
													1328	=>X"00",
													1329	=>X"00",
													1330	=>X"00",
													1331	=>X"00",
													1332	=>X"00",
													1333	=>X"00",
													1334	=>X"00",
													1335	=>X"00",
													1336	=>X"00",
													1337	=>X"00",
													1338	=>X"00",
													1339	=>X"00",
													1340	=>X"00",
													1341	=>X"00",
													1342	=>X"00",
													1343	=>X"00",
													1344	=>X"00",
													1345	=>X"00",
													1346	=>X"00",
													1347	=>X"00",
													1348	=>X"00",
													1349	=>X"00",
													1350	=>X"00",
													1351	=>X"00",
													1352	=>X"00",
													1353	=>X"00",
													1354	=>X"00",
													1355	=>X"00",
													1356	=>X"00",
													1357	=>X"00",
													1358	=>X"00",
													1359	=>X"00",
													1360	=>X"00",
													1361	=>X"00",
													1362	=>X"00",
													1363	=>X"00",
													1364	=>X"00",
													1365	=>X"00",
													1366	=>X"00",
													1367	=>X"00",
													1368	=>X"00",
													1369	=>X"00",
													1370	=>X"00",
													1371	=>X"00",
													1372	=>X"00",
													1373	=>X"00",
													1374	=>X"00",
													1375	=>X"00",
													1376	=>X"00",
													1377	=>X"00",
													1378	=>X"00",
													1379	=>X"00",
													1380	=>X"00",
													1381	=>X"00",
													1382	=>X"00",
													1383	=>X"00",
													1384	=>X"00",
													1385	=>X"00",
													1386	=>X"00",
													1387	=>X"00",
													1388	=>X"00",
													1389	=>X"00",
													1390	=>X"00",
													1391	=>X"00",
													1392	=>X"00",
													1393	=>X"00",
													1394	=>X"00",
													1395	=>X"00",
													1396	=>X"00",
													1397	=>X"00",
													1398	=>X"00",
													1399	=>X"00",
													1400	=>X"00",
													1401	=>X"00",
													1402	=>X"00",
													1403	=>X"00",
													1404	=>X"00",
													1405	=>X"00",
													1406	=>X"00",
													1407	=>X"00",
													1408	=>X"00",
													1409	=>X"00",
													1410	=>X"00",
													1411	=>X"00",
													1412	=>X"00",
													1413	=>X"00",
													1414	=>X"00",
													1415	=>X"00",
													1416	=>X"00",
													1417	=>X"00",
													1418	=>X"00",
													1419	=>X"00",
													1420	=>X"00",
													1421	=>X"00",
													1422	=>X"00",
													1423	=>X"00",
													1424	=>X"00",
													1425	=>X"00",
													1426	=>X"00",
													1427	=>X"00",
													1428	=>X"00",
													1429	=>X"00",
													1430	=>X"00",
													1431	=>X"00",
													1432	=>X"00",
													1433	=>X"00",
													1434	=>X"00",
													1435	=>X"00",
													1436	=>X"00",
													1437	=>X"00",
													1438	=>X"00",
													1439	=>X"00",
													1440	=>X"00",
													1441	=>X"00",
													1442	=>X"00",
													1443	=>X"00",
													1444	=>X"00",
													1445	=>X"00",
													1446	=>X"00",
													1447	=>X"00",
													1448	=>X"00",
													1449	=>X"00",
													1450	=>X"00",
													1451	=>X"00",
													1452	=>X"00",
													1453	=>X"00",
													1454	=>X"00",
													1455	=>X"00",
													1456	=>X"00",
													1457	=>X"00",
													1458	=>X"00",
													1459	=>X"00",
													1460	=>X"00",
													1461	=>X"00",
													1462	=>X"00",
													1463	=>X"00",
													1464	=>X"00",
													1465	=>X"00",
													1466	=>X"00",
													1467	=>X"00",
													1468	=>X"00",
													1469	=>X"00",
													1470	=>X"00",
													1471	=>X"00",
													1472	=>X"00",
													1473	=>X"00",
													1474	=>X"00",
													1475	=>X"00",
													1476	=>X"00",
													1477	=>X"00",
													1478	=>X"00",
													1479	=>X"00",
													1480	=>X"00",
													1481	=>X"00",
													1482	=>X"00",
													1483	=>X"00",
													1484	=>X"00",
													1485	=>X"00",
													1486	=>X"00",
													1487	=>X"00",
													1488	=>X"00",
													1489	=>X"00",
													1490	=>X"00",
													1491	=>X"00",
													1492	=>X"00",
													1493	=>X"00",
													1494	=>X"00",
													1495	=>X"00",
													1496	=>X"00",
													1497	=>X"00",
													1498	=>X"00",
													1499	=>X"00",
													1500	=>X"00",
													1501	=>X"00",
													1502	=>X"00",
													1503	=>X"00",
													1504	=>X"00",
													1505	=>X"00",
													1506	=>X"00",
													1507	=>X"00",
													1508	=>X"00",
													1509	=>X"00",
													1510	=>X"00",
													1511	=>X"00",
													1512	=>X"00",
													1513	=>X"00",
													1514	=>X"00",
													1515	=>X"00",
													1516	=>X"00",
													1517	=>X"00",
													1518	=>X"00",
													1519	=>X"00",
													1520	=>X"00",
													1521	=>X"00",
													1522	=>X"00",
													1523	=>X"00",
													1524	=>X"00",
													1525	=>X"00",
													1526	=>X"00",
													1527	=>X"00",
													1528	=>X"00",
													1529	=>X"00",
													1530	=>X"00",
													1531	=>X"00",
													1532	=>X"00",
													1533	=>X"00",
													1534	=>X"00",
													1535	=>X"00",
													1536	=>X"00",
													1537	=>X"00",
													1538	=>X"00",
													1539	=>X"00",
													1540	=>X"00",
													1541	=>X"00",
													1542	=>X"00",
													1543	=>X"00",
													1544	=>X"00",
													1545	=>X"00",
													1546	=>X"00",
													1547	=>X"00",
													1548	=>X"00",
													1549	=>X"00",
													1550	=>X"00",
													1551	=>X"00",
													1552	=>X"00",
													1553	=>X"00",
													1554	=>X"00",
													1555	=>X"00",
													1556	=>X"00",
													1557	=>X"00",
													1558	=>X"00",
													1559	=>X"00",
													1560	=>X"00",
													1561	=>X"00",
													1562	=>X"00",
													1563	=>X"00",
													1564	=>X"00",
													1565	=>X"00",
													1566	=>X"00",
													1567	=>X"00",
													1568	=>X"00",
													1569	=>X"00",
													1570	=>X"00",
													1571	=>X"00",
													1572	=>X"00",
													1573	=>X"00",
													1574	=>X"00",
													1575	=>X"00",
													1576	=>X"00",
													1577	=>X"00",
													1578	=>X"00",
													1579	=>X"00",
													1580	=>X"00",
													1581	=>X"00",
													1582	=>X"00",
													1583	=>X"00",
													1584	=>X"00",
													1585	=>X"00",
													1586	=>X"00",
													1587	=>X"00",
													1588	=>X"00",
													1589	=>X"00",
													1590	=>X"00",
													1591	=>X"00",
													1592	=>X"00",
													1593	=>X"00",
													1594	=>X"00",
													1595	=>X"00",
													1596	=>X"00",
													1597	=>X"00",
													1598	=>X"00",
													1599	=>X"00",
													1600	=>X"00",
													1601	=>X"00",
													1602	=>X"00",
													1603	=>X"00",
													1604	=>X"00",
													1605	=>X"00",
													1606	=>X"00",
													1607	=>X"00",
													1608	=>X"00",
													1609	=>X"00",
													1610	=>X"00",
													1611	=>X"00",
													1612	=>X"00",
													1613	=>X"00",
													1614	=>X"00",
													1615	=>X"00",
													1616	=>X"00",
													1617	=>X"00",
													1618	=>X"00",
													1619	=>X"00",
													1620	=>X"00",
													1621	=>X"00",
													1622	=>X"00",
													1623	=>X"00",
													1624	=>X"00",
													1625	=>X"00",
													1626	=>X"00",
													1627	=>X"00",
													1628	=>X"00",
													1629	=>X"00",
													1630	=>X"00",
													1631	=>X"07",
													1632	=>X"ff",
													1633	=>X"f8",
													1634	=>X"00",
													1635	=>X"00",
													1636	=>X"00",
													1637	=>X"00",
													1638	=>X"00",
													1639	=>X"00",
													1640	=>X"00",
													1641	=>X"00",
													1642	=>X"00",
													1643	=>X"00",
													1644	=>X"00",
													1645	=>X"00",
													1646	=>X"00",
													1647	=>X"00",
													1648	=>X"00",
													1649	=>X"00",
													1650	=>X"00",
													1651	=>X"00",
													1652	=>X"00",
													1653	=>X"00",
													1654	=>X"00",
													1655	=>X"00",
													1656	=>X"00",
													1657	=>X"00",
													1658	=>X"00",
													1659	=>X"00",
													1660	=>X"00",
													1661	=>X"00",
													1662	=>X"00",
													1663	=>X"00",
													1664	=>X"00",
													1665	=>X"00",
													1666	=>X"00",
													1667	=>X"00",
													1668	=>X"00",
													1669	=>X"00",
													1670	=>X"00",
													1671	=>X"0f",
													1672	=>X"ff",
													1673	=>X"fc",
													1674	=>X"00",
													1675	=>X"00",
													1676	=>X"00",
													1677	=>X"00",
													1678	=>X"00",
													1679	=>X"00",
													1680	=>X"00",
													1681	=>X"00",
													1682	=>X"00",
													1683	=>X"00",
													1684	=>X"00",
													1685	=>X"00",
													1686	=>X"00",
													1687	=>X"00",
													1688	=>X"00",
													1689	=>X"00",
													1690	=>X"00",
													1691	=>X"00",
													1692	=>X"00",
													1693	=>X"00",
													1694	=>X"00",
													1695	=>X"00",
													1696	=>X"00",
													1697	=>X"00",
													1698	=>X"00",
													1699	=>X"00",
													1700	=>X"00",
													1701	=>X"00",
													1702	=>X"00",
													1703	=>X"00",
													1704	=>X"00",
													1705	=>X"00",
													1706	=>X"00",
													1707	=>X"00",
													1708	=>X"00",
													1709	=>X"00",
													1710	=>X"00",
													1711	=>X"1f",
													1712	=>X"ff",
													1713	=>X"fe",
													1714	=>X"00",
													1715	=>X"00",
													1716	=>X"00",
													1717	=>X"00",
													1718	=>X"00",
													1719	=>X"00",
													1720	=>X"00",
													1721	=>X"00",
													1722	=>X"00",
													1723	=>X"00",
													1724	=>X"00",
													1725	=>X"00",
													1726	=>X"00",
													1727	=>X"00",
													1728	=>X"00",
													1729	=>X"00",
													1730	=>X"00",
													1731	=>X"00",
													1732	=>X"00",
													1733	=>X"00",
													1734	=>X"00",
													1735	=>X"00",
													1736	=>X"00",
													1737	=>X"00",
													1738	=>X"00",
													1739	=>X"00",
													1740	=>X"00",
													1741	=>X"00",
													1742	=>X"00",
													1743	=>X"00",
													1744	=>X"00",
													1745	=>X"00",
													1746	=>X"00",
													1747	=>X"00",
													1748	=>X"00",
													1749	=>X"00",
													1750	=>X"00",
													1751	=>X"1f",
													1752	=>X"ff",
													1753	=>X"fe",
													1754	=>X"00",
													1755	=>X"00",
													1756	=>X"00",
													1757	=>X"00",
													1758	=>X"00",
													1759	=>X"00",
													1760	=>X"00",
													1761	=>X"00",
													1762	=>X"00",
													1763	=>X"00",
													1764	=>X"00",
													1765	=>X"00",
													1766	=>X"00",
													1767	=>X"00",
													1768	=>X"00",
													1769	=>X"00",
													1770	=>X"00",
													1771	=>X"00",
													1772	=>X"00",
													1773	=>X"00",
													1774	=>X"00",
													1775	=>X"00",
													1776	=>X"00",
													1777	=>X"00",
													1778	=>X"00",
													1779	=>X"00",
													1780	=>X"00",
													1781	=>X"00",
													1782	=>X"00",
													1783	=>X"00",
													1784	=>X"00",
													1785	=>X"00",
													1786	=>X"00",
													1787	=>X"00",
													1788	=>X"00",
													1789	=>X"00",
													1790	=>X"00",
													1791	=>X"3f",
													1792	=>X"ff",
													1793	=>X"ff",
													1794	=>X"00",
													1795	=>X"00",
													1796	=>X"00",
													1797	=>X"00",
													1798	=>X"00",
													1799	=>X"00",
													1800	=>X"00",
													1801	=>X"00",
													1802	=>X"00",
													1803	=>X"00",
													1804	=>X"00",
													1805	=>X"00",
													1806	=>X"00",
													1807	=>X"00",
													1808	=>X"00",
													1809	=>X"00",
													1810	=>X"00",
													1811	=>X"00",
													1812	=>X"00",
													1813	=>X"00",
													1814	=>X"00",
													1815	=>X"00",
													1816	=>X"00",
													1817	=>X"00",
													1818	=>X"00",
													1819	=>X"00",
													1820	=>X"00",
													1821	=>X"00",
													1822	=>X"00",
													1823	=>X"00",
													1824	=>X"00",
													1825	=>X"00",
													1826	=>X"00",
													1827	=>X"00",
													1828	=>X"00",
													1829	=>X"00",
													1830	=>X"00",
													1831	=>X"7f",
													1832	=>X"ff",
													1833	=>X"ff",
													1834	=>X"80",
													1835	=>X"00",
													1836	=>X"00",
													1837	=>X"00",
													1838	=>X"00",
													1839	=>X"00",
													1840	=>X"00",
													1841	=>X"00",
													1842	=>X"00",
													1843	=>X"00",
													1844	=>X"00",
													1845	=>X"00",
													1846	=>X"00",
													1847	=>X"00",
													1848	=>X"00",
													1849	=>X"00",
													1850	=>X"00",
													1851	=>X"00",
													1852	=>X"00",
													1853	=>X"00",
													1854	=>X"00",
													1855	=>X"00",
													1856	=>X"00",
													1857	=>X"00",
													1858	=>X"00",
													1859	=>X"00",
													1860	=>X"00",
													1861	=>X"00",
													1862	=>X"00",
													1863	=>X"00",
													1864	=>X"00",
													1865	=>X"00",
													1866	=>X"00",
													1867	=>X"00",
													1868	=>X"00",
													1869	=>X"00",
													1870	=>X"00",
													1871	=>X"7f",
													1872	=>X"ff",
													1873	=>X"ff",
													1874	=>X"80",
													1875	=>X"00",
													1876	=>X"00",
													1877	=>X"00",
													1878	=>X"00",
													1879	=>X"00",
													1880	=>X"00",
													1881	=>X"00",
													1882	=>X"00",
													1883	=>X"00",
													1884	=>X"00",
													1885	=>X"00",
													1886	=>X"00",
													1887	=>X"00",
													1888	=>X"00",
													1889	=>X"00",
													1890	=>X"00",
													1891	=>X"00",
													1892	=>X"00",
													1893	=>X"00",
													1894	=>X"00",
													1895	=>X"00",
													1896	=>X"00",
													1897	=>X"00",
													1898	=>X"00",
													1899	=>X"00",
													1900	=>X"00",
													1901	=>X"00",
													1902	=>X"00",
													1903	=>X"00",
													1904	=>X"00",
													1905	=>X"00",
													1906	=>X"00",
													1907	=>X"00",
													1908	=>X"00",
													1909	=>X"00",
													1910	=>X"00",
													1911	=>X"ff",
													1912	=>X"ff",
													1913	=>X"ff",
													1914	=>X"c0",
													1915	=>X"00",
													1916	=>X"00",
													1917	=>X"00",
													1918	=>X"00",
													1919	=>X"00",
													1920	=>X"00",
													1921	=>X"00",
													1922	=>X"00",
													1923	=>X"00",
													1924	=>X"00",
													1925	=>X"00",
													1926	=>X"00",
													1927	=>X"00",
													1928	=>X"00",
													1929	=>X"00",
													1930	=>X"00",
													1931	=>X"00",
													1932	=>X"00",
													1933	=>X"00",
													1934	=>X"00",
													1935	=>X"00",
													1936	=>X"00",
													1937	=>X"00",
													1938	=>X"00",
													1939	=>X"00",
													1940	=>X"00",
													1941	=>X"00",
													1942	=>X"00",
													1943	=>X"00",
													1944	=>X"00",
													1945	=>X"00",
													1946	=>X"00",
													1947	=>X"00",
													1948	=>X"00",
													1949	=>X"00",
													1950	=>X"00",
													1951	=>X"ff",
													1952	=>X"ff",
													1953	=>X"ff",
													1954	=>X"c0",
													1955	=>X"00",
													1956	=>X"00",
													1957	=>X"00",
													1958	=>X"00",
													1959	=>X"00",
													1960	=>X"00",
													1961	=>X"00",
													1962	=>X"00",
													1963	=>X"00",
													1964	=>X"00",
													1965	=>X"00",
													1966	=>X"00",
													1967	=>X"00",
													1968	=>X"00",
													1969	=>X"00",
													1970	=>X"00",
													1971	=>X"00",
													1972	=>X"00",
													1973	=>X"00",
													1974	=>X"00",
													1975	=>X"00",
													1976	=>X"00",
													1977	=>X"00",
													1978	=>X"00",
													1979	=>X"00",
													1980	=>X"00",
													1981	=>X"00",
													1982	=>X"00",
													1983	=>X"00",
													1984	=>X"00",
													1985	=>X"00",
													1986	=>X"00",
													1987	=>X"00",
													1988	=>X"00",
													1989	=>X"00",
													1990	=>X"01",
													1991	=>X"fc",
													1992	=>X"00",
													1993	=>X"1f",
													1994	=>X"e0",
													1995	=>X"00",
													1996	=>X"00",
													1997	=>X"00",
													1998	=>X"00",
													1999	=>X"00",
													2000	=>X"00",
													2001	=>X"00",
													2002	=>X"00",
													2003	=>X"00",
													2004	=>X"00",
													2005	=>X"00",
													2006	=>X"00",
													2007	=>X"00",
													2008	=>X"00",
													2009	=>X"00",
													2010	=>X"00",
													2011	=>X"00",
													2012	=>X"00",
													2013	=>X"00",
													2014	=>X"00",
													2015	=>X"00",
													2016	=>X"00",
													2017	=>X"00",
													2018	=>X"00",
													2019	=>X"00",
													2020	=>X"00",
													2021	=>X"00",
													2022	=>X"00",
													2023	=>X"00",
													2024	=>X"00",
													2025	=>X"00",
													2026	=>X"00",
													2027	=>X"00",
													2028	=>X"00",
													2029	=>X"00",
													2030	=>X"01",
													2031	=>X"f8",
													2032	=>X"f8",
													2033	=>X"0f",
													2034	=>X"e0",
													2035	=>X"00",
													2036	=>X"00",
													2037	=>X"00",
													2038	=>X"00",
													2039	=>X"00",
													2040	=>X"00",
													2041	=>X"00",
													2042	=>X"00",
													2043	=>X"00",
													2044	=>X"00",
													2045	=>X"00",
													2046	=>X"00",
													2047	=>X"00",
													2048	=>X"00",
													2049	=>X"00",
													2050	=>X"00",
													2051	=>X"00",
													2052	=>X"00",
													2053	=>X"00",
													2054	=>X"00",
													2055	=>X"00",
													2056	=>X"00",
													2057	=>X"00",
													2058	=>X"00",
													2059	=>X"00",
													2060	=>X"00",
													2061	=>X"00",
													2062	=>X"00",
													2063	=>X"00",
													2064	=>X"00",
													2065	=>X"00",
													2066	=>X"00",
													2067	=>X"00",
													2068	=>X"00",
													2069	=>X"00",
													2070	=>X"03",
													2071	=>X"f9",
													2072	=>X"f0",
													2073	=>X"07",
													2074	=>X"f0",
													2075	=>X"00",
													2076	=>X"00",
													2077	=>X"00",
													2078	=>X"00",
													2079	=>X"00",
													2080	=>X"00",
													2081	=>X"00",
													2082	=>X"00",
													2083	=>X"00",
													2084	=>X"00",
													2085	=>X"00",
													2086	=>X"00",
													2087	=>X"00",
													2088	=>X"00",
													2089	=>X"00",
													2090	=>X"00",
													2091	=>X"00",
													2092	=>X"00",
													2093	=>X"00",
													2094	=>X"00",
													2095	=>X"00",
													2096	=>X"00",
													2097	=>X"00",
													2098	=>X"00",
													2099	=>X"00",
													2100	=>X"00",
													2101	=>X"00",
													2102	=>X"00",
													2103	=>X"00",
													2104	=>X"00",
													2105	=>X"00",
													2106	=>X"00",
													2107	=>X"00",
													2108	=>X"00",
													2109	=>X"00",
													2110	=>X"03",
													2111	=>X"f3",
													2112	=>X"e0",
													2113	=>X"c7",
													2114	=>X"f0",
													2115	=>X"00",
													2116	=>X"00",
													2117	=>X"00",
													2118	=>X"00",
													2119	=>X"00",
													2120	=>X"00",
													2121	=>X"00",
													2122	=>X"00",
													2123	=>X"00",
													2124	=>X"00",
													2125	=>X"00",
													2126	=>X"00",
													2127	=>X"00",
													2128	=>X"00",
													2129	=>X"00",
													2130	=>X"00",
													2131	=>X"00",
													2132	=>X"00",
													2133	=>X"00",
													2134	=>X"00",
													2135	=>X"00",
													2136	=>X"00",
													2137	=>X"00",
													2138	=>X"00",
													2139	=>X"00",
													2140	=>X"00",
													2141	=>X"00",
													2142	=>X"00",
													2143	=>X"00",
													2144	=>X"00",
													2145	=>X"00",
													2146	=>X"00",
													2147	=>X"00",
													2148	=>X"00",
													2149	=>X"00",
													2150	=>X"07",
													2151	=>X"e3",
													2152	=>X"c0",
													2153	=>X"f3",
													2154	=>X"f0",
													2155	=>X"00",
													2156	=>X"00",
													2157	=>X"00",
													2158	=>X"00",
													2159	=>X"00",
													2160	=>X"00",
													2161	=>X"00",
													2162	=>X"00",
													2163	=>X"00",
													2164	=>X"00",
													2165	=>X"00",
													2166	=>X"00",
													2167	=>X"00",
													2168	=>X"00",
													2169	=>X"00",
													2170	=>X"00",
													2171	=>X"00",
													2172	=>X"00",
													2173	=>X"00",
													2174	=>X"00",
													2175	=>X"00",
													2176	=>X"00",
													2177	=>X"00",
													2178	=>X"00",
													2179	=>X"00",
													2180	=>X"00",
													2181	=>X"00",
													2182	=>X"00",
													2183	=>X"00",
													2184	=>X"00",
													2185	=>X"00",
													2186	=>X"00",
													2187	=>X"00",
													2188	=>X"00",
													2189	=>X"00",
													2190	=>X"07",
													2191	=>X"e7",
													2192	=>X"80",
													2193	=>X"7b",
													2194	=>X"f8",
													2195	=>X"00",
													2196	=>X"00",
													2197	=>X"00",
													2198	=>X"00",
													2199	=>X"00",
													2200	=>X"00",
													2201	=>X"00",
													2202	=>X"00",
													2203	=>X"00",
													2204	=>X"00",
													2205	=>X"00",
													2206	=>X"00",
													2207	=>X"00",
													2208	=>X"00",
													2209	=>X"00",
													2210	=>X"00",
													2211	=>X"00",
													2212	=>X"00",
													2213	=>X"00",
													2214	=>X"00",
													2215	=>X"00",
													2216	=>X"00",
													2217	=>X"00",
													2218	=>X"00",
													2219	=>X"00",
													2220	=>X"00",
													2221	=>X"00",
													2222	=>X"00",
													2223	=>X"00",
													2224	=>X"00",
													2225	=>X"00",
													2226	=>X"00",
													2227	=>X"00",
													2228	=>X"00",
													2229	=>X"00",
													2230	=>X"07",
													2231	=>X"c7",
													2232	=>X"80",
													2233	=>X"39",
													2234	=>X"f8",
													2235	=>X"00",
													2236	=>X"00",
													2237	=>X"00",
													2238	=>X"00",
													2239	=>X"00",
													2240	=>X"00",
													2241	=>X"00",
													2242	=>X"00",
													2243	=>X"00",
													2244	=>X"00",
													2245	=>X"00",
													2246	=>X"00",
													2247	=>X"00",
													2248	=>X"00",
													2249	=>X"00",
													2250	=>X"00",
													2251	=>X"00",
													2252	=>X"00",
													2253	=>X"00",
													2254	=>X"00",
													2255	=>X"00",
													2256	=>X"00",
													2257	=>X"00",
													2258	=>X"00",
													2259	=>X"00",
													2260	=>X"00",
													2261	=>X"00",
													2262	=>X"00",
													2263	=>X"00",
													2264	=>X"00",
													2265	=>X"00",
													2266	=>X"00",
													2267	=>X"00",
													2268	=>X"00",
													2269	=>X"00",
													2270	=>X"0f",
													2271	=>X"c7",
													2272	=>X"07",
													2273	=>X"1d",
													2274	=>X"fc",
													2275	=>X"00",
													2276	=>X"00",
													2277	=>X"00",
													2278	=>X"00",
													2279	=>X"00",
													2280	=>X"00",
													2281	=>X"00",
													2282	=>X"00",
													2283	=>X"00",
													2284	=>X"00",
													2285	=>X"00",
													2286	=>X"00",
													2287	=>X"00",
													2288	=>X"00",
													2289	=>X"00",
													2290	=>X"00",
													2291	=>X"00",
													2292	=>X"00",
													2293	=>X"00",
													2294	=>X"00",
													2295	=>X"00",
													2296	=>X"00",
													2297	=>X"00",
													2298	=>X"00",
													2299	=>X"00",
													2300	=>X"00",
													2301	=>X"00",
													2302	=>X"00",
													2303	=>X"00",
													2304	=>X"00",
													2305	=>X"00",
													2306	=>X"00",
													2307	=>X"00",
													2308	=>X"00",
													2309	=>X"00",
													2310	=>X"0f",
													2311	=>X"c7",
													2312	=>X"07",
													2313	=>X"1c",
													2314	=>X"fc",
													2315	=>X"00",
													2316	=>X"00",
													2317	=>X"00",
													2318	=>X"00",
													2319	=>X"00",
													2320	=>X"00",
													2321	=>X"00",
													2322	=>X"00",
													2323	=>X"00",
													2324	=>X"00",
													2325	=>X"00",
													2326	=>X"00",
													2327	=>X"00",
													2328	=>X"00",
													2329	=>X"00",
													2330	=>X"00",
													2331	=>X"00",
													2332	=>X"00",
													2333	=>X"00",
													2334	=>X"00",
													2335	=>X"00",
													2336	=>X"00",
													2337	=>X"00",
													2338	=>X"00",
													2339	=>X"00",
													2340	=>X"00",
													2341	=>X"00",
													2342	=>X"00",
													2343	=>X"00",
													2344	=>X"00",
													2345	=>X"00",
													2346	=>X"00",
													2347	=>X"00",
													2348	=>X"00",
													2349	=>X"00",
													2350	=>X"1f",
													2351	=>X"8e",
													2352	=>X"07",
													2353	=>X"1e",
													2354	=>X"fc",
													2355	=>X"00",
													2356	=>X"00",
													2357	=>X"00",
													2358	=>X"00",
													2359	=>X"00",
													2360	=>X"00",
													2361	=>X"00",
													2362	=>X"00",
													2363	=>X"00",
													2364	=>X"00",
													2365	=>X"00",
													2366	=>X"00",
													2367	=>X"00",
													2368	=>X"00",
													2369	=>X"00",
													2370	=>X"00",
													2371	=>X"00",
													2372	=>X"00",
													2373	=>X"00",
													2374	=>X"00",
													2375	=>X"00",
													2376	=>X"00",
													2377	=>X"00",
													2378	=>X"00",
													2379	=>X"00",
													2380	=>X"00",
													2381	=>X"00",
													2382	=>X"00",
													2383	=>X"00",
													2384	=>X"00",
													2385	=>X"00",
													2386	=>X"00",
													2387	=>X"00",
													2388	=>X"00",
													2389	=>X"00",
													2390	=>X"1f",
													2391	=>X"8e",
													2392	=>X"07",
													2393	=>X"0e",
													2394	=>X"7e",
													2395	=>X"00",
													2396	=>X"00",
													2397	=>X"00",
													2398	=>X"00",
													2399	=>X"00",
													2400	=>X"00",
													2401	=>X"00",
													2402	=>X"00",
													2403	=>X"00",
													2404	=>X"00",
													2405	=>X"00",
													2406	=>X"00",
													2407	=>X"00",
													2408	=>X"00",
													2409	=>X"00",
													2410	=>X"00",
													2411	=>X"00",
													2412	=>X"00",
													2413	=>X"00",
													2414	=>X"00",
													2415	=>X"00",
													2416	=>X"00",
													2417	=>X"00",
													2418	=>X"00",
													2419	=>X"00",
													2420	=>X"00",
													2421	=>X"00",
													2422	=>X"00",
													2423	=>X"00",
													2424	=>X"00",
													2425	=>X"00",
													2426	=>X"00",
													2427	=>X"00",
													2428	=>X"00",
													2429	=>X"00",
													2430	=>X"1f",
													2431	=>X"0e",
													2432	=>X"07",
													2433	=>X"0e",
													2434	=>X"7e",
													2435	=>X"00",
													2436	=>X"00",
													2437	=>X"00",
													2438	=>X"00",
													2439	=>X"00",
													2440	=>X"00",
													2441	=>X"00",
													2442	=>X"00",
													2443	=>X"00",
													2444	=>X"00",
													2445	=>X"00",
													2446	=>X"00",
													2447	=>X"00",
													2448	=>X"00",
													2449	=>X"00",
													2450	=>X"00",
													2451	=>X"00",
													2452	=>X"00",
													2453	=>X"00",
													2454	=>X"00",
													2455	=>X"00",
													2456	=>X"00",
													2457	=>X"00",
													2458	=>X"00",
													2459	=>X"00",
													2460	=>X"00",
													2461	=>X"00",
													2462	=>X"00",
													2463	=>X"00",
													2464	=>X"00",
													2465	=>X"00",
													2466	=>X"00",
													2467	=>X"00",
													2468	=>X"00",
													2469	=>X"00",
													2470	=>X"1f",
													2471	=>X"0f",
													2472	=>X"07",
													2473	=>X"0e",
													2474	=>X"7e",
													2475	=>X"00",
													2476	=>X"00",
													2477	=>X"00",
													2478	=>X"00",
													2479	=>X"00",
													2480	=>X"00",
													2481	=>X"00",
													2482	=>X"00",
													2483	=>X"00",
													2484	=>X"00",
													2485	=>X"00",
													2486	=>X"00",
													2487	=>X"00",
													2488	=>X"00",
													2489	=>X"00",
													2490	=>X"00",
													2491	=>X"00",
													2492	=>X"00",
													2493	=>X"00",
													2494	=>X"00",
													2495	=>X"00",
													2496	=>X"00",
													2497	=>X"00",
													2498	=>X"00",
													2499	=>X"00",
													2500	=>X"00",
													2501	=>X"00",
													2502	=>X"00",
													2503	=>X"00",
													2504	=>X"00",
													2505	=>X"00",
													2506	=>X"00",
													2507	=>X"00",
													2508	=>X"00",
													2509	=>X"00",
													2510	=>X"3f",
													2511	=>X"0f",
													2512	=>X"07",
													2513	=>X"0e",
													2514	=>X"3e",
													2515	=>X"00",
													2516	=>X"00",
													2517	=>X"00",
													2518	=>X"00",
													2519	=>X"00",
													2520	=>X"00",
													2521	=>X"00",
													2522	=>X"00",
													2523	=>X"00",
													2524	=>X"00",
													2525	=>X"00",
													2526	=>X"00",
													2527	=>X"00",
													2528	=>X"00",
													2529	=>X"00",
													2530	=>X"00",
													2531	=>X"00",
													2532	=>X"00",
													2533	=>X"00",
													2534	=>X"00",
													2535	=>X"00",
													2536	=>X"00",
													2537	=>X"00",
													2538	=>X"00",
													2539	=>X"00",
													2540	=>X"00",
													2541	=>X"00",
													2542	=>X"00",
													2543	=>X"00",
													2544	=>X"00",
													2545	=>X"00",
													2546	=>X"00",
													2547	=>X"00",
													2548	=>X"00",
													2549	=>X"00",
													2550	=>X"3e",
													2551	=>X"0f",
													2552	=>X"07",
													2553	=>X"0e",
													2554	=>X"3f",
													2555	=>X"00",
													2556	=>X"00",
													2557	=>X"00",
													2558	=>X"00",
													2559	=>X"00",
													2560	=>X"00",
													2561	=>X"00",
													2562	=>X"00",
													2563	=>X"00",
													2564	=>X"00",
													2565	=>X"00",
													2566	=>X"00",
													2567	=>X"00",
													2568	=>X"00",
													2569	=>X"00",
													2570	=>X"00",
													2571	=>X"00",
													2572	=>X"00",
													2573	=>X"00",
													2574	=>X"00",
													2575	=>X"00",
													2576	=>X"00",
													2577	=>X"00",
													2578	=>X"00",
													2579	=>X"00",
													2580	=>X"00",
													2581	=>X"00",
													2582	=>X"00",
													2583	=>X"00",
													2584	=>X"00",
													2585	=>X"00",
													2586	=>X"00",
													2587	=>X"00",
													2588	=>X"00",
													2589	=>X"00",
													2590	=>X"3e",
													2591	=>X"07",
													2592	=>X"e7",
													2593	=>X"1e",
													2594	=>X"3f",
													2595	=>X"00",
													2596	=>X"00",
													2597	=>X"00",
													2598	=>X"00",
													2599	=>X"00",
													2600	=>X"00",
													2601	=>X"00",
													2602	=>X"00",
													2603	=>X"00",
													2604	=>X"00",
													2605	=>X"00",
													2606	=>X"00",
													2607	=>X"00",
													2608	=>X"00",
													2609	=>X"00",
													2610	=>X"00",
													2611	=>X"00",
													2612	=>X"00",
													2613	=>X"00",
													2614	=>X"00",
													2615	=>X"00",
													2616	=>X"00",
													2617	=>X"00",
													2618	=>X"00",
													2619	=>X"00",
													2620	=>X"00",
													2621	=>X"00",
													2622	=>X"00",
													2623	=>X"00",
													2624	=>X"00",
													2625	=>X"00",
													2626	=>X"00",
													2627	=>X"00",
													2628	=>X"00",
													2629	=>X"00",
													2630	=>X"7e",
													2631	=>X"07",
													2632	=>X"ff",
													2633	=>X"7e",
													2634	=>X"1f",
													2635	=>X"00",
													2636	=>X"00",
													2637	=>X"00",
													2638	=>X"00",
													2639	=>X"00",
													2640	=>X"00",
													2641	=>X"00",
													2642	=>X"00",
													2643	=>X"00",
													2644	=>X"00",
													2645	=>X"00",
													2646	=>X"00",
													2647	=>X"00",
													2648	=>X"00",
													2649	=>X"00",
													2650	=>X"00",
													2651	=>X"00",
													2652	=>X"00",
													2653	=>X"00",
													2654	=>X"00",
													2655	=>X"00",
													2656	=>X"00",
													2657	=>X"00",
													2658	=>X"00",
													2659	=>X"00",
													2660	=>X"00",
													2661	=>X"00",
													2662	=>X"00",
													2663	=>X"00",
													2664	=>X"00",
													2665	=>X"00",
													2666	=>X"00",
													2667	=>X"00",
													2668	=>X"00",
													2669	=>X"00",
													2670	=>X"7e",
													2671	=>X"07",
													2672	=>X"ff",
													2673	=>X"fe",
													2674	=>X"1f",
													2675	=>X"80",
													2676	=>X"00",
													2677	=>X"00",
													2678	=>X"00",
													2679	=>X"00",
													2680	=>X"00",
													2681	=>X"00",
													2682	=>X"00",
													2683	=>X"00",
													2684	=>X"00",
													2685	=>X"00",
													2686	=>X"00",
													2687	=>X"00",
													2688	=>X"00",
													2689	=>X"00",
													2690	=>X"00",
													2691	=>X"00",
													2692	=>X"00",
													2693	=>X"00",
													2694	=>X"00",
													2695	=>X"00",
													2696	=>X"00",
													2697	=>X"00",
													2698	=>X"00",
													2699	=>X"00",
													2700	=>X"00",
													2701	=>X"00",
													2702	=>X"00",
													2703	=>X"00",
													2704	=>X"00",
													2705	=>X"00",
													2706	=>X"00",
													2707	=>X"00",
													2708	=>X"00",
													2709	=>X"00",
													2710	=>X"7c",
													2711	=>X"03",
													2712	=>X"ff",
													2713	=>X"fe",
													2714	=>X"1f",
													2715	=>X"80",
													2716	=>X"00",
													2717	=>X"00",
													2718	=>X"00",
													2719	=>X"00",
													2720	=>X"00",
													2721	=>X"00",
													2722	=>X"00",
													2723	=>X"00",
													2724	=>X"00",
													2725	=>X"00",
													2726	=>X"00",
													2727	=>X"00",
													2728	=>X"00",
													2729	=>X"00",
													2730	=>X"00",
													2731	=>X"00",
													2732	=>X"00",
													2733	=>X"00",
													2734	=>X"00",
													2735	=>X"00",
													2736	=>X"00",
													2737	=>X"00",
													2738	=>X"00",
													2739	=>X"00",
													2740	=>X"00",
													2741	=>X"00",
													2742	=>X"00",
													2743	=>X"00",
													2744	=>X"00",
													2745	=>X"00",
													2746	=>X"00",
													2747	=>X"00",
													2748	=>X"00",
													2749	=>X"00",
													2750	=>X"7c",
													2751	=>X"01",
													2752	=>X"ff",
													2753	=>X"fc",
													2754	=>X"1f",
													2755	=>X"80",
													2756	=>X"00",
													2757	=>X"00",
													2758	=>X"00",
													2759	=>X"00",
													2760	=>X"00",
													2761	=>X"00",
													2762	=>X"00",
													2763	=>X"00",
													2764	=>X"00",
													2765	=>X"00",
													2766	=>X"00",
													2767	=>X"00",
													2768	=>X"00",
													2769	=>X"00",
													2770	=>X"00",
													2771	=>X"00",
													2772	=>X"00",
													2773	=>X"00",
													2774	=>X"00",
													2775	=>X"00",
													2776	=>X"00",
													2777	=>X"00",
													2778	=>X"00",
													2779	=>X"00",
													2780	=>X"00",
													2781	=>X"00",
													2782	=>X"00",
													2783	=>X"00",
													2784	=>X"00",
													2785	=>X"00",
													2786	=>X"00",
													2787	=>X"00",
													2788	=>X"00",
													2789	=>X"00",
													2790	=>X"fc",
													2791	=>X"00",
													2792	=>X"7f",
													2793	=>X"fc",
													2794	=>X"0f",
													2795	=>X"80",
													2796	=>X"00",
													2797	=>X"00",
													2798	=>X"00",
													2799	=>X"00",
													2800	=>X"00",
													2801	=>X"00",
													2802	=>X"00",
													2803	=>X"00",
													2804	=>X"00",
													2805	=>X"00",
													2806	=>X"00",
													2807	=>X"00",
													2808	=>X"00",
													2809	=>X"00",
													2810	=>X"00",
													2811	=>X"00",
													2812	=>X"00",
													2813	=>X"00",
													2814	=>X"00",
													2815	=>X"00",
													2816	=>X"00",
													2817	=>X"00",
													2818	=>X"00",
													2819	=>X"00",
													2820	=>X"00",
													2821	=>X"00",
													2822	=>X"00",
													2823	=>X"00",
													2824	=>X"00",
													2825	=>X"00",
													2826	=>X"00",
													2827	=>X"00",
													2828	=>X"00",
													2829	=>X"00",
													2830	=>X"fc",
													2831	=>X"00",
													2832	=>X"1f",
													2833	=>X"f0",
													2834	=>X"0f",
													2835	=>X"80",
													2836	=>X"00",
													2837	=>X"00",
													2838	=>X"00",
													2839	=>X"00",
													2840	=>X"00",
													2841	=>X"00",
													2842	=>X"00",
													2843	=>X"00",
													2844	=>X"00",
													2845	=>X"00",
													2846	=>X"00",
													2847	=>X"00",
													2848	=>X"00",
													2849	=>X"00",
													2850	=>X"00",
													2851	=>X"00",
													2852	=>X"00",
													2853	=>X"00",
													2854	=>X"00",
													2855	=>X"00",
													2856	=>X"00",
													2857	=>X"00",
													2858	=>X"00",
													2859	=>X"00",
													2860	=>X"00",
													2861	=>X"00",
													2862	=>X"00",
													2863	=>X"00",
													2864	=>X"00",
													2865	=>X"00",
													2866	=>X"00",
													2867	=>X"00",
													2868	=>X"00",
													2869	=>X"00",
													2870	=>X"f8",
													2871	=>X"7c",
													2872	=>X"00",
													2873	=>X"80",
													2874	=>X"0f",
													2875	=>X"c0",
													2876	=>X"00",
													2877	=>X"00",
													2878	=>X"00",
													2879	=>X"00",
													2880	=>X"00",
													2881	=>X"00",
													2882	=>X"00",
													2883	=>X"00",
													2884	=>X"00",
													2885	=>X"00",
													2886	=>X"00",
													2887	=>X"00",
													2888	=>X"00",
													2889	=>X"00",
													2890	=>X"00",
													2891	=>X"00",
													2892	=>X"00",
													2893	=>X"00",
													2894	=>X"00",
													2895	=>X"00",
													2896	=>X"00",
													2897	=>X"00",
													2898	=>X"00",
													2899	=>X"00",
													2900	=>X"00",
													2901	=>X"00",
													2902	=>X"00",
													2903	=>X"00",
													2904	=>X"00",
													2905	=>X"00",
													2906	=>X"00",
													2907	=>X"00",
													2908	=>X"00",
													2909	=>X"00",
													2910	=>X"f8",
													2911	=>X"7f",
													2912	=>X"80",
													2913	=>X"00",
													2914	=>X"0f",
													2915	=>X"c0",
													2916	=>X"00",
													2917	=>X"00",
													2918	=>X"00",
													2919	=>X"00",
													2920	=>X"00",
													2921	=>X"00",
													2922	=>X"00",
													2923	=>X"00",
													2924	=>X"00",
													2925	=>X"00",
													2926	=>X"00",
													2927	=>X"00",
													2928	=>X"00",
													2929	=>X"00",
													2930	=>X"00",
													2931	=>X"00",
													2932	=>X"00",
													2933	=>X"00",
													2934	=>X"00",
													2935	=>X"00",
													2936	=>X"00",
													2937	=>X"00",
													2938	=>X"00",
													2939	=>X"00",
													2940	=>X"00",
													2941	=>X"00",
													2942	=>X"00",
													2943	=>X"00",
													2944	=>X"00",
													2945	=>X"00",
													2946	=>X"00",
													2947	=>X"00",
													2948	=>X"00",
													2949	=>X"00",
													2950	=>X"f8",
													2951	=>X"7f",
													2952	=>X"f0",
													2953	=>X"00",
													2954	=>X"07",
													2955	=>X"c0",
													2956	=>X"00",
													2957	=>X"00",
													2958	=>X"00",
													2959	=>X"00",
													2960	=>X"00",
													2961	=>X"00",
													2962	=>X"00",
													2963	=>X"00",
													2964	=>X"00",
													2965	=>X"00",
													2966	=>X"00",
													2967	=>X"00",
													2968	=>X"00",
													2969	=>X"00",
													2970	=>X"00",
													2971	=>X"00",
													2972	=>X"00",
													2973	=>X"00",
													2974	=>X"00",
													2975	=>X"00",
													2976	=>X"00",
													2977	=>X"00",
													2978	=>X"00",
													2979	=>X"00",
													2980	=>X"00",
													2981	=>X"00",
													2982	=>X"00",
													2983	=>X"00",
													2984	=>X"00",
													2985	=>X"00",
													2986	=>X"00",
													2987	=>X"00",
													2988	=>X"00",
													2989	=>X"01",
													2990	=>X"f8",
													2991	=>X"ff",
													2992	=>X"fc",
													2993	=>X"00",
													2994	=>X"07",
													2995	=>X"c0",
													2996	=>X"00",
													2997	=>X"00",
													2998	=>X"00",
													2999	=>X"00",
													3000	=>X"00",
													3001	=>X"00",
													3002	=>X"00",
													3003	=>X"00",
													3004	=>X"00",
													3005	=>X"00",
													3006	=>X"00",
													3007	=>X"00",
													3008	=>X"00",
													3009	=>X"00",
													3010	=>X"00",
													3011	=>X"00",
													3012	=>X"00",
													3013	=>X"00",
													3014	=>X"00",
													3015	=>X"00",
													3016	=>X"00",
													3017	=>X"00",
													3018	=>X"00",
													3019	=>X"00",
													3020	=>X"00",
													3021	=>X"00",
													3022	=>X"00",
													3023	=>X"00",
													3024	=>X"00",
													3025	=>X"00",
													3026	=>X"00",
													3027	=>X"00",
													3028	=>X"00",
													3029	=>X"01",
													3030	=>X"f0",
													3031	=>X"ff",
													3032	=>X"ff",
													3033	=>X"00",
													3034	=>X"07",
													3035	=>X"c0",
													3036	=>X"00",
													3037	=>X"00",
													3038	=>X"00",
													3039	=>X"00",
													3040	=>X"00",
													3041	=>X"00",
													3042	=>X"00",
													3043	=>X"00",
													3044	=>X"00",
													3045	=>X"00",
													3046	=>X"00",
													3047	=>X"00",
													3048	=>X"00",
													3049	=>X"00",
													3050	=>X"00",
													3051	=>X"00",
													3052	=>X"00",
													3053	=>X"00",
													3054	=>X"00",
													3055	=>X"00",
													3056	=>X"00",
													3057	=>X"00",
													3058	=>X"00",
													3059	=>X"00",
													3060	=>X"00",
													3061	=>X"00",
													3062	=>X"00",
													3063	=>X"00",
													3064	=>X"00",
													3065	=>X"00",
													3066	=>X"00",
													3067	=>X"00",
													3068	=>X"00",
													3069	=>X"01",
													3070	=>X"f0",
													3071	=>X"c0",
													3072	=>X"7f",
													3073	=>X"c0",
													3074	=>X"07",
													3075	=>X"e0",
													3076	=>X"00",
													3077	=>X"00",
													3078	=>X"00",
													3079	=>X"00",
													3080	=>X"00",
													3081	=>X"00",
													3082	=>X"00",
													3083	=>X"00",
													3084	=>X"00",
													3085	=>X"00",
													3086	=>X"00",
													3087	=>X"00",
													3088	=>X"00",
													3089	=>X"00",
													3090	=>X"00",
													3091	=>X"00",
													3092	=>X"00",
													3093	=>X"00",
													3094	=>X"00",
													3095	=>X"00",
													3096	=>X"00",
													3097	=>X"00",
													3098	=>X"00",
													3099	=>X"00",
													3100	=>X"00",
													3101	=>X"00",
													3102	=>X"00",
													3103	=>X"00",
													3104	=>X"00",
													3105	=>X"00",
													3106	=>X"00",
													3107	=>X"00",
													3108	=>X"00",
													3109	=>X"01",
													3110	=>X"f0",
													3111	=>X"00",
													3112	=>X"0f",
													3113	=>X"e0",
													3114	=>X"07",
													3115	=>X"e0",
													3116	=>X"00",
													3117	=>X"00",
													3118	=>X"00",
													3119	=>X"00",
													3120	=>X"00",
													3121	=>X"00",
													3122	=>X"00",
													3123	=>X"00",
													3124	=>X"00",
													3125	=>X"00",
													3126	=>X"00",
													3127	=>X"00",
													3128	=>X"00",
													3129	=>X"00",
													3130	=>X"00",
													3131	=>X"00",
													3132	=>X"00",
													3133	=>X"00",
													3134	=>X"00",
													3135	=>X"00",
													3136	=>X"00",
													3137	=>X"00",
													3138	=>X"00",
													3139	=>X"00",
													3140	=>X"00",
													3141	=>X"00",
													3142	=>X"00",
													3143	=>X"00",
													3144	=>X"00",
													3145	=>X"00",
													3146	=>X"00",
													3147	=>X"00",
													3148	=>X"00",
													3149	=>X"01",
													3150	=>X"f0",
													3151	=>X"00",
													3152	=>X"03",
													3153	=>X"f8",
													3154	=>X"03",
													3155	=>X"e0",
													3156	=>X"00",
													3157	=>X"00",
													3158	=>X"00",
													3159	=>X"00",
													3160	=>X"00",
													3161	=>X"00",
													3162	=>X"00",
													3163	=>X"00",
													3164	=>X"00",
													3165	=>X"00",
													3166	=>X"00",
													3167	=>X"00",
													3168	=>X"00",
													3169	=>X"00",
													3170	=>X"00",
													3171	=>X"00",
													3172	=>X"00",
													3173	=>X"00",
													3174	=>X"00",
													3175	=>X"00",
													3176	=>X"00",
													3177	=>X"00",
													3178	=>X"00",
													3179	=>X"00",
													3180	=>X"00",
													3181	=>X"00",
													3182	=>X"00",
													3183	=>X"00",
													3184	=>X"00",
													3185	=>X"00",
													3186	=>X"00",
													3187	=>X"00",
													3188	=>X"00",
													3189	=>X"03",
													3190	=>X"f0",
													3191	=>X"00",
													3192	=>X"01",
													3193	=>X"fc",
													3194	=>X"03",
													3195	=>X"e0",
													3196	=>X"00",
													3197	=>X"00",
													3198	=>X"00",
													3199	=>X"00",
													3200	=>X"00",
													3201	=>X"00",
													3202	=>X"00",
													3203	=>X"00",
													3204	=>X"00",
													3205	=>X"00",
													3206	=>X"00",
													3207	=>X"00",
													3208	=>X"00",
													3209	=>X"00",
													3210	=>X"00",
													3211	=>X"00",
													3212	=>X"00",
													3213	=>X"00",
													3214	=>X"00",
													3215	=>X"00",
													3216	=>X"00",
													3217	=>X"00",
													3218	=>X"00",
													3219	=>X"00",
													3220	=>X"00",
													3221	=>X"00",
													3222	=>X"00",
													3223	=>X"00",
													3224	=>X"00",
													3225	=>X"00",
													3226	=>X"00",
													3227	=>X"00",
													3228	=>X"00",
													3229	=>X"03",
													3230	=>X"e0",
													3231	=>X"00",
													3232	=>X"00",
													3233	=>X"7e",
													3234	=>X"43",
													3235	=>X"e0",
													3236	=>X"00",
													3237	=>X"00",
													3238	=>X"00",
													3239	=>X"00",
													3240	=>X"00",
													3241	=>X"00",
													3242	=>X"00",
													3243	=>X"00",
													3244	=>X"00",
													3245	=>X"00",
													3246	=>X"00",
													3247	=>X"00",
													3248	=>X"00",
													3249	=>X"00",
													3250	=>X"00",
													3251	=>X"00",
													3252	=>X"00",
													3253	=>X"00",
													3254	=>X"00",
													3255	=>X"00",
													3256	=>X"00",
													3257	=>X"00",
													3258	=>X"00",
													3259	=>X"00",
													3260	=>X"00",
													3261	=>X"00",
													3262	=>X"00",
													3263	=>X"00",
													3264	=>X"00",
													3265	=>X"00",
													3266	=>X"00",
													3267	=>X"00",
													3268	=>X"00",
													3269	=>X"03",
													3270	=>X"e0",
													3271	=>X"80",
													3272	=>X"00",
													3273	=>X"1f",
													3274	=>X"e3",
													3275	=>X"e0",
													3276	=>X"00",
													3277	=>X"00",
													3278	=>X"00",
													3279	=>X"00",
													3280	=>X"00",
													3281	=>X"00",
													3282	=>X"00",
													3283	=>X"00",
													3284	=>X"00",
													3285	=>X"00",
													3286	=>X"00",
													3287	=>X"00",
													3288	=>X"00",
													3289	=>X"00",
													3290	=>X"00",
													3291	=>X"00",
													3292	=>X"00",
													3293	=>X"00",
													3294	=>X"00",
													3295	=>X"00",
													3296	=>X"00",
													3297	=>X"00",
													3298	=>X"00",
													3299	=>X"00",
													3300	=>X"00",
													3301	=>X"00",
													3302	=>X"00",
													3303	=>X"00",
													3304	=>X"00",
													3305	=>X"00",
													3306	=>X"00",
													3307	=>X"00",
													3308	=>X"00",
													3309	=>X"03",
													3310	=>X"e1",
													3311	=>X"80",
													3312	=>X"00",
													3313	=>X"0f",
													3314	=>X"e3",
													3315	=>X"f0",
													3316	=>X"00",
													3317	=>X"00",
													3318	=>X"00",
													3319	=>X"00",
													3320	=>X"00",
													3321	=>X"00",
													3322	=>X"00",
													3323	=>X"00",
													3324	=>X"00",
													3325	=>X"00",
													3326	=>X"00",
													3327	=>X"00",
													3328	=>X"00",
													3329	=>X"00",
													3330	=>X"00",
													3331	=>X"00",
													3332	=>X"00",
													3333	=>X"00",
													3334	=>X"00",
													3335	=>X"00",
													3336	=>X"00",
													3337	=>X"00",
													3338	=>X"00",
													3339	=>X"00",
													3340	=>X"00",
													3341	=>X"00",
													3342	=>X"00",
													3343	=>X"00",
													3344	=>X"00",
													3345	=>X"00",
													3346	=>X"00",
													3347	=>X"00",
													3348	=>X"00",
													3349	=>X"03",
													3350	=>X"e1",
													3351	=>X"e0",
													3352	=>X"00",
													3353	=>X"07",
													3354	=>X"e3",
													3355	=>X"f0",
													3356	=>X"00",
													3357	=>X"00",
													3358	=>X"00",
													3359	=>X"00",
													3360	=>X"00",
													3361	=>X"00",
													3362	=>X"00",
													3363	=>X"00",
													3364	=>X"00",
													3365	=>X"00",
													3366	=>X"00",
													3367	=>X"00",
													3368	=>X"00",
													3369	=>X"00",
													3370	=>X"00",
													3371	=>X"00",
													3372	=>X"00",
													3373	=>X"00",
													3374	=>X"00",
													3375	=>X"00",
													3376	=>X"00",
													3377	=>X"00",
													3378	=>X"00",
													3379	=>X"00",
													3380	=>X"00",
													3381	=>X"00",
													3382	=>X"00",
													3383	=>X"00",
													3384	=>X"00",
													3385	=>X"00",
													3386	=>X"00",
													3387	=>X"00",
													3388	=>X"00",
													3389	=>X"03",
													3390	=>X"e1",
													3391	=>X"fc",
													3392	=>X"00",
													3393	=>X"01",
													3394	=>X"e3",
													3395	=>X"f0",
													3396	=>X"00",
													3397	=>X"00",
													3398	=>X"00",
													3399	=>X"00",
													3400	=>X"00",
													3401	=>X"00",
													3402	=>X"00",
													3403	=>X"00",
													3404	=>X"00",
													3405	=>X"00",
													3406	=>X"00",
													3407	=>X"00",
													3408	=>X"00",
													3409	=>X"00",
													3410	=>X"00",
													3411	=>X"00",
													3412	=>X"00",
													3413	=>X"00",
													3414	=>X"00",
													3415	=>X"00",
													3416	=>X"00",
													3417	=>X"00",
													3418	=>X"00",
													3419	=>X"00",
													3420	=>X"00",
													3421	=>X"00",
													3422	=>X"00",
													3423	=>X"00",
													3424	=>X"00",
													3425	=>X"00",
													3426	=>X"00",
													3427	=>X"00",
													3428	=>X"00",
													3429	=>X"07",
													3430	=>X"e1",
													3431	=>X"ff",
													3432	=>X"c0",
													3433	=>X"01",
													3434	=>X"e1",
													3435	=>X"f0",
													3436	=>X"00",
													3437	=>X"00",
													3438	=>X"00",
													3439	=>X"00",
													3440	=>X"00",
													3441	=>X"00",
													3442	=>X"00",
													3443	=>X"00",
													3444	=>X"00",
													3445	=>X"00",
													3446	=>X"00",
													3447	=>X"00",
													3448	=>X"00",
													3449	=>X"00",
													3450	=>X"00",
													3451	=>X"00",
													3452	=>X"00",
													3453	=>X"00",
													3454	=>X"00",
													3455	=>X"00",
													3456	=>X"00",
													3457	=>X"00",
													3458	=>X"00",
													3459	=>X"00",
													3460	=>X"00",
													3461	=>X"00",
													3462	=>X"00",
													3463	=>X"00",
													3464	=>X"00",
													3465	=>X"00",
													3466	=>X"00",
													3467	=>X"00",
													3468	=>X"00",
													3469	=>X"07",
													3470	=>X"e1",
													3471	=>X"ff",
													3472	=>X"fe",
													3473	=>X"01",
													3474	=>X"e1",
													3475	=>X"f0",
													3476	=>X"00",
													3477	=>X"00",
													3478	=>X"00",
													3479	=>X"00",
													3480	=>X"00",
													3481	=>X"00",
													3482	=>X"00",
													3483	=>X"00",
													3484	=>X"00",
													3485	=>X"00",
													3486	=>X"00",
													3487	=>X"00",
													3488	=>X"00",
													3489	=>X"00",
													3490	=>X"00",
													3491	=>X"00",
													3492	=>X"00",
													3493	=>X"00",
													3494	=>X"00",
													3495	=>X"00",
													3496	=>X"00",
													3497	=>X"00",
													3498	=>X"00",
													3499	=>X"00",
													3500	=>X"00",
													3501	=>X"00",
													3502	=>X"00",
													3503	=>X"00",
													3504	=>X"00",
													3505	=>X"00",
													3506	=>X"00",
													3507	=>X"00",
													3508	=>X"00",
													3509	=>X"07",
													3510	=>X"c1",
													3511	=>X"ff",
													3512	=>X"ff",
													3513	=>X"f1",
													3514	=>X"e1",
													3515	=>X"f0",
													3516	=>X"00",
													3517	=>X"00",
													3518	=>X"00",
													3519	=>X"00",
													3520	=>X"00",
													3521	=>X"00",
													3522	=>X"00",
													3523	=>X"00",
													3524	=>X"00",
													3525	=>X"00",
													3526	=>X"00",
													3527	=>X"00",
													3528	=>X"00",
													3529	=>X"00",
													3530	=>X"00",
													3531	=>X"00",
													3532	=>X"00",
													3533	=>X"00",
													3534	=>X"00",
													3535	=>X"00",
													3536	=>X"00",
													3537	=>X"00",
													3538	=>X"00",
													3539	=>X"00",
													3540	=>X"00",
													3541	=>X"00",
													3542	=>X"00",
													3543	=>X"00",
													3544	=>X"00",
													3545	=>X"00",
													3546	=>X"00",
													3547	=>X"00",
													3548	=>X"00",
													3549	=>X"07",
													3550	=>X"c1",
													3551	=>X"bf",
													3552	=>X"ff",
													3553	=>X"ff",
													3554	=>X"e1",
													3555	=>X"f0",
													3556	=>X"00",
													3557	=>X"00",
													3558	=>X"00",
													3559	=>X"00",
													3560	=>X"00",
													3561	=>X"00",
													3562	=>X"00",
													3563	=>X"00",
													3564	=>X"00",
													3565	=>X"00",
													3566	=>X"00",
													3567	=>X"00",
													3568	=>X"00",
													3569	=>X"00",
													3570	=>X"00",
													3571	=>X"00",
													3572	=>X"00",
													3573	=>X"00",
													3574	=>X"00",
													3575	=>X"00",
													3576	=>X"00",
													3577	=>X"00",
													3578	=>X"00",
													3579	=>X"00",
													3580	=>X"00",
													3581	=>X"00",
													3582	=>X"00",
													3583	=>X"00",
													3584	=>X"00",
													3585	=>X"00",
													3586	=>X"00",
													3587	=>X"00",
													3588	=>X"00",
													3589	=>X"07",
													3590	=>X"c1",
													3591	=>X"83",
													3592	=>X"ff",
													3593	=>X"ff",
													3594	=>X"e1",
													3595	=>X"f8",
													3596	=>X"00",
													3597	=>X"00",
													3598	=>X"00",
													3599	=>X"00",
													3600	=>X"00",
													3601	=>X"00",
													3602	=>X"00",
													3603	=>X"00",
													3604	=>X"00",
													3605	=>X"00",
													3606	=>X"00",
													3607	=>X"00",
													3608	=>X"00",
													3609	=>X"00",
													3610	=>X"00",
													3611	=>X"00",
													3612	=>X"00",
													3613	=>X"00",
													3614	=>X"00",
													3615	=>X"00",
													3616	=>X"00",
													3617	=>X"00",
													3618	=>X"00",
													3619	=>X"00",
													3620	=>X"00",
													3621	=>X"00",
													3622	=>X"00",
													3623	=>X"00",
													3624	=>X"00",
													3625	=>X"00",
													3626	=>X"00",
													3627	=>X"00",
													3628	=>X"00",
													3629	=>X"07",
													3630	=>X"c0",
													3631	=>X"00",
													3632	=>X"1f",
													3633	=>X"ff",
													3634	=>X"e1",
													3635	=>X"f8",
													3636	=>X"00",
													3637	=>X"00",
													3638	=>X"00",
													3639	=>X"00",
													3640	=>X"00",
													3641	=>X"00",
													3642	=>X"00",
													3643	=>X"00",
													3644	=>X"00",
													3645	=>X"00",
													3646	=>X"00",
													3647	=>X"00",
													3648	=>X"00",
													3649	=>X"00",
													3650	=>X"00",
													3651	=>X"00",
													3652	=>X"00",
													3653	=>X"00",
													3654	=>X"00",
													3655	=>X"00",
													3656	=>X"00",
													3657	=>X"00",
													3658	=>X"00",
													3659	=>X"00",
													3660	=>X"00",
													3661	=>X"00",
													3662	=>X"00",
													3663	=>X"00",
													3664	=>X"00",
													3665	=>X"00",
													3666	=>X"00",
													3667	=>X"00",
													3668	=>X"00",
													3669	=>X"07",
													3670	=>X"c0",
													3671	=>X"00",
													3672	=>X"01",
													3673	=>X"ff",
													3674	=>X"e1",
													3675	=>X"f8",
													3676	=>X"00",
													3677	=>X"00",
													3678	=>X"00",
													3679	=>X"00",
													3680	=>X"00",
													3681	=>X"00",
													3682	=>X"00",
													3683	=>X"00",
													3684	=>X"00",
													3685	=>X"00",
													3686	=>X"00",
													3687	=>X"00",
													3688	=>X"00",
													3689	=>X"00",
													3690	=>X"00",
													3691	=>X"00",
													3692	=>X"00",
													3693	=>X"00",
													3694	=>X"00",
													3695	=>X"00",
													3696	=>X"00",
													3697	=>X"00",
													3698	=>X"00",
													3699	=>X"00",
													3700	=>X"00",
													3701	=>X"00",
													3702	=>X"00",
													3703	=>X"00",
													3704	=>X"00",
													3705	=>X"00",
													3706	=>X"00",
													3707	=>X"00",
													3708	=>X"00",
													3709	=>X"07",
													3710	=>X"c0",
													3711	=>X"00",
													3712	=>X"00",
													3713	=>X"1f",
													3714	=>X"e1",
													3715	=>X"f8",
													3716	=>X"00",
													3717	=>X"00",
													3718	=>X"00",
													3719	=>X"00",
													3720	=>X"00",
													3721	=>X"00",
													3722	=>X"00",
													3723	=>X"00",
													3724	=>X"00",
													3725	=>X"00",
													3726	=>X"00",
													3727	=>X"00",
													3728	=>X"00",
													3729	=>X"00",
													3730	=>X"00",
													3731	=>X"00",
													3732	=>X"00",
													3733	=>X"00",
													3734	=>X"00",
													3735	=>X"00",
													3736	=>X"00",
													3737	=>X"00",
													3738	=>X"00",
													3739	=>X"00",
													3740	=>X"00",
													3741	=>X"00",
													3742	=>X"00",
													3743	=>X"00",
													3744	=>X"00",
													3745	=>X"00",
													3746	=>X"00",
													3747	=>X"00",
													3748	=>X"00",
													3749	=>X"07",
													3750	=>X"c0",
													3751	=>X"00",
													3752	=>X"00",
													3753	=>X"00",
													3754	=>X"e0",
													3755	=>X"f8",
													3756	=>X"00",
													3757	=>X"00",
													3758	=>X"00",
													3759	=>X"00",
													3760	=>X"00",
													3761	=>X"00",
													3762	=>X"00",
													3763	=>X"00",
													3764	=>X"00",
													3765	=>X"00",
													3766	=>X"00",
													3767	=>X"00",
													3768	=>X"00",
													3769	=>X"00",
													3770	=>X"00",
													3771	=>X"00",
													3772	=>X"00",
													3773	=>X"00",
													3774	=>X"00",
													3775	=>X"00",
													3776	=>X"00",
													3777	=>X"00",
													3778	=>X"00",
													3779	=>X"00",
													3780	=>X"00",
													3781	=>X"00",
													3782	=>X"00",
													3783	=>X"00",
													3784	=>X"00",
													3785	=>X"00",
													3786	=>X"00",
													3787	=>X"00",
													3788	=>X"00",
													3789	=>X"0f",
													3790	=>X"c0",
													3791	=>X"00",
													3792	=>X"00",
													3793	=>X"00",
													3794	=>X"60",
													3795	=>X"f8",
													3796	=>X"00",
													3797	=>X"00",
													3798	=>X"00",
													3799	=>X"00",
													3800	=>X"00",
													3801	=>X"00",
													3802	=>X"00",
													3803	=>X"00",
													3804	=>X"00",
													3805	=>X"00",
													3806	=>X"00",
													3807	=>X"00",
													3808	=>X"00",
													3809	=>X"00",
													3810	=>X"00",
													3811	=>X"00",
													3812	=>X"00",
													3813	=>X"00",
													3814	=>X"00",
													3815	=>X"00",
													3816	=>X"00",
													3817	=>X"00",
													3818	=>X"00",
													3819	=>X"00",
													3820	=>X"00",
													3821	=>X"00",
													3822	=>X"00",
													3823	=>X"00",
													3824	=>X"00",
													3825	=>X"00",
													3826	=>X"00",
													3827	=>X"00",
													3828	=>X"00",
													3829	=>X"0f",
													3830	=>X"c0",
													3831	=>X"0f",
													3832	=>X"ff",
													3833	=>X"00",
													3834	=>X"60",
													3835	=>X"f8",
													3836	=>X"00",
													3837	=>X"00",
													3838	=>X"00",
													3839	=>X"00",
													3840	=>X"00",
													3841	=>X"00",
													3842	=>X"00",
													3843	=>X"00",
													3844	=>X"00",
													3845	=>X"00",
													3846	=>X"00",
													3847	=>X"00",
													3848	=>X"00",
													3849	=>X"00",
													3850	=>X"00",
													3851	=>X"00",
													3852	=>X"00",
													3853	=>X"00",
													3854	=>X"00",
													3855	=>X"00",
													3856	=>X"00",
													3857	=>X"00",
													3858	=>X"00",
													3859	=>X"00",
													3860	=>X"00",
													3861	=>X"00",
													3862	=>X"00",
													3863	=>X"00",
													3864	=>X"00",
													3865	=>X"00",
													3866	=>X"00",
													3867	=>X"00",
													3868	=>X"00",
													3869	=>X"0f",
													3870	=>X"80",
													3871	=>X"3f",
													3872	=>X"ff",
													3873	=>X"e0",
													3874	=>X"00",
													3875	=>X"f8",
													3876	=>X"00",
													3877	=>X"00",
													3878	=>X"00",
													3879	=>X"00",
													3880	=>X"00",
													3881	=>X"00",
													3882	=>X"00",
													3883	=>X"00",
													3884	=>X"00",
													3885	=>X"00",
													3886	=>X"00",
													3887	=>X"00",
													3888	=>X"00",
													3889	=>X"00",
													3890	=>X"00",
													3891	=>X"00",
													3892	=>X"00",
													3893	=>X"00",
													3894	=>X"00",
													3895	=>X"00",
													3896	=>X"00",
													3897	=>X"00",
													3898	=>X"00",
													3899	=>X"00",
													3900	=>X"00",
													3901	=>X"00",
													3902	=>X"00",
													3903	=>X"00",
													3904	=>X"00",
													3905	=>X"00",
													3906	=>X"00",
													3907	=>X"00",
													3908	=>X"00",
													3909	=>X"0f",
													3910	=>X"80",
													3911	=>X"ff",
													3912	=>X"ff",
													3913	=>X"f8",
													3914	=>X"00",
													3915	=>X"f8",
													3916	=>X"00",
													3917	=>X"00",
													3918	=>X"00",
													3919	=>X"00",
													3920	=>X"00",
													3921	=>X"00",
													3922	=>X"00",
													3923	=>X"00",
													3924	=>X"00",
													3925	=>X"00",
													3926	=>X"00",
													3927	=>X"00",
													3928	=>X"00",
													3929	=>X"00",
													3930	=>X"00",
													3931	=>X"00",
													3932	=>X"00",
													3933	=>X"00",
													3934	=>X"00",
													3935	=>X"00",
													3936	=>X"00",
													3937	=>X"00",
													3938	=>X"00",
													3939	=>X"00",
													3940	=>X"00",
													3941	=>X"00",
													3942	=>X"00",
													3943	=>X"00",
													3944	=>X"00",
													3945	=>X"00",
													3946	=>X"00",
													3947	=>X"00",
													3948	=>X"00",
													3949	=>X"0f",
													3950	=>X"80",
													3951	=>X"ff",
													3952	=>X"ff",
													3953	=>X"fe",
													3954	=>X"00",
													3955	=>X"f8",
													3956	=>X"00",
													3957	=>X"00",
													3958	=>X"00",
													3959	=>X"00",
													3960	=>X"00",
													3961	=>X"00",
													3962	=>X"00",
													3963	=>X"00",
													3964	=>X"00",
													3965	=>X"00",
													3966	=>X"00",
													3967	=>X"00",
													3968	=>X"00",
													3969	=>X"00",
													3970	=>X"00",
													3971	=>X"00",
													3972	=>X"00",
													3973	=>X"00",
													3974	=>X"00",
													3975	=>X"00",
													3976	=>X"00",
													3977	=>X"00",
													3978	=>X"00",
													3979	=>X"00",
													3980	=>X"00",
													3981	=>X"00",
													3982	=>X"00",
													3983	=>X"00",
													3984	=>X"00",
													3985	=>X"00",
													3986	=>X"00",
													3987	=>X"00",
													3988	=>X"00",
													3989	=>X"0f",
													3990	=>X"81",
													3991	=>X"ff",
													3992	=>X"ff",
													3993	=>X"ff",
													3994	=>X"00",
													3995	=>X"f8",
													3996	=>X"00",
													3997	=>X"00",
													3998	=>X"00",
													3999	=>X"00",
													4000	=>X"00",
													4001	=>X"00",
													4002	=>X"00",
													4003	=>X"00",
													4004	=>X"00",
													4005	=>X"00",
													4006	=>X"00",
													4007	=>X"00",
													4008	=>X"00",
													4009	=>X"00",
													4010	=>X"00",
													4011	=>X"00",
													4012	=>X"00",
													4013	=>X"00",
													4014	=>X"00",
													4015	=>X"00",
													4016	=>X"00",
													4017	=>X"00",
													4018	=>X"00",
													4019	=>X"00",
													4020	=>X"00",
													4021	=>X"00",
													4022	=>X"00",
													4023	=>X"00",
													4024	=>X"00",
													4025	=>X"00",
													4026	=>X"00",
													4027	=>X"00",
													4028	=>X"00",
													4029	=>X"0f",
													4030	=>X"81",
													4031	=>X"fe",
													4032	=>X"03",
													4033	=>X"ff",
													4034	=>X"80",
													4035	=>X"f8",
													4036	=>X"00",
													4037	=>X"00",
													4038	=>X"00",
													4039	=>X"00",
													4040	=>X"00",
													4041	=>X"00",
													4042	=>X"00",
													4043	=>X"00",
													4044	=>X"00",
													4045	=>X"00",
													4046	=>X"00",
													4047	=>X"00",
													4048	=>X"00",
													4049	=>X"00",
													4050	=>X"00",
													4051	=>X"00",
													4052	=>X"00",
													4053	=>X"00",
													4054	=>X"00",
													4055	=>X"00",
													4056	=>X"00",
													4057	=>X"00",
													4058	=>X"00",
													4059	=>X"00",
													4060	=>X"00",
													4061	=>X"00",
													4062	=>X"00",
													4063	=>X"00",
													4064	=>X"00",
													4065	=>X"00",
													4066	=>X"00",
													4067	=>X"00",
													4068	=>X"00",
													4069	=>X"0f",
													4070	=>X"83",
													4071	=>X"f0",
													4072	=>X"00",
													4073	=>X"7f",
													4074	=>X"80",
													4075	=>X"fc",
													4076	=>X"00",
													4077	=>X"00",
													4078	=>X"00",
													4079	=>X"00",
													4080	=>X"00",
													4081	=>X"00",
													4082	=>X"00",
													4083	=>X"00",
													4084	=>X"00",
													4085	=>X"00",
													4086	=>X"00",
													4087	=>X"00",
													4088	=>X"00",
													4089	=>X"00",
													4090	=>X"00",
													4091	=>X"00",
													4092	=>X"00",
													4093	=>X"00",
													4094	=>X"00",
													4095	=>X"00",
													4096	=>X"00",
													4097	=>X"00",
													4098	=>X"00",
													4099	=>X"00",
													4100	=>X"00",
													4101	=>X"00",
													4102	=>X"00",
													4103	=>X"00",
													4104	=>X"00",
													4105	=>X"00",
													4106	=>X"00",
													4107	=>X"00",
													4108	=>X"00",
													4109	=>X"0f",
													4110	=>X"83",
													4111	=>X"e0",
													4112	=>X"00",
													4113	=>X"1f",
													4114	=>X"c0",
													4115	=>X"fc",
													4116	=>X"00",
													4117	=>X"00",
													4118	=>X"00",
													4119	=>X"00",
													4120	=>X"00",
													4121	=>X"00",
													4122	=>X"00",
													4123	=>X"00",
													4124	=>X"00",
													4125	=>X"00",
													4126	=>X"00",
													4127	=>X"00",
													4128	=>X"00",
													4129	=>X"00",
													4130	=>X"00",
													4131	=>X"00",
													4132	=>X"00",
													4133	=>X"00",
													4134	=>X"00",
													4135	=>X"00",
													4136	=>X"00",
													4137	=>X"00",
													4138	=>X"00",
													4139	=>X"00",
													4140	=>X"00",
													4141	=>X"00",
													4142	=>X"00",
													4143	=>X"00",
													4144	=>X"00",
													4145	=>X"00",
													4146	=>X"00",
													4147	=>X"00",
													4148	=>X"00",
													4149	=>X"0f",
													4150	=>X"83",
													4151	=>X"c0",
													4152	=>X"00",
													4153	=>X"0f",
													4154	=>X"e0",
													4155	=>X"fc",
													4156	=>X"00",
													4157	=>X"00",
													4158	=>X"00",
													4159	=>X"00",
													4160	=>X"00",
													4161	=>X"00",
													4162	=>X"00",
													4163	=>X"00",
													4164	=>X"00",
													4165	=>X"00",
													4166	=>X"00",
													4167	=>X"00",
													4168	=>X"00",
													4169	=>X"00",
													4170	=>X"00",
													4171	=>X"00",
													4172	=>X"00",
													4173	=>X"00",
													4174	=>X"00",
													4175	=>X"00",
													4176	=>X"00",
													4177	=>X"00",
													4178	=>X"00",
													4179	=>X"00",
													4180	=>X"00",
													4181	=>X"00",
													4182	=>X"00",
													4183	=>X"00",
													4184	=>X"00",
													4185	=>X"00",
													4186	=>X"00",
													4187	=>X"00",
													4188	=>X"00",
													4189	=>X"1f",
													4190	=>X"83",
													4191	=>X"c0",
													4192	=>X"00",
													4193	=>X"03",
													4194	=>X"e0",
													4195	=>X"fc",
													4196	=>X"00",
													4197	=>X"00",
													4198	=>X"00",
													4199	=>X"00",
													4200	=>X"00",
													4201	=>X"00",
													4202	=>X"00",
													4203	=>X"00",
													4204	=>X"00",
													4205	=>X"00",
													4206	=>X"00",
													4207	=>X"00",
													4208	=>X"00",
													4209	=>X"00",
													4210	=>X"00",
													4211	=>X"00",
													4212	=>X"00",
													4213	=>X"00",
													4214	=>X"00",
													4215	=>X"00",
													4216	=>X"00",
													4217	=>X"00",
													4218	=>X"00",
													4219	=>X"00",
													4220	=>X"00",
													4221	=>X"00",
													4222	=>X"00",
													4223	=>X"00",
													4224	=>X"00",
													4225	=>X"00",
													4226	=>X"00",
													4227	=>X"00",
													4228	=>X"00",
													4229	=>X"1f",
													4230	=>X"83",
													4231	=>X"c0",
													4232	=>X"00",
													4233	=>X"01",
													4234	=>X"e0",
													4235	=>X"fc",
													4236	=>X"00",
													4237	=>X"00",
													4238	=>X"00",
													4239	=>X"00",
													4240	=>X"00",
													4241	=>X"00",
													4242	=>X"00",
													4243	=>X"00",
													4244	=>X"00",
													4245	=>X"00",
													4246	=>X"00",
													4247	=>X"00",
													4248	=>X"00",
													4249	=>X"00",
													4250	=>X"00",
													4251	=>X"00",
													4252	=>X"00",
													4253	=>X"00",
													4254	=>X"00",
													4255	=>X"00",
													4256	=>X"00",
													4257	=>X"00",
													4258	=>X"00",
													4259	=>X"00",
													4260	=>X"00",
													4261	=>X"00",
													4262	=>X"00",
													4263	=>X"00",
													4264	=>X"00",
													4265	=>X"00",
													4266	=>X"00",
													4267	=>X"00",
													4268	=>X"00",
													4269	=>X"1f",
													4270	=>X"83",
													4271	=>X"c0",
													4272	=>X"00",
													4273	=>X"01",
													4274	=>X"e0",
													4275	=>X"fc",
													4276	=>X"00",
													4277	=>X"00",
													4278	=>X"00",
													4279	=>X"00",
													4280	=>X"00",
													4281	=>X"00",
													4282	=>X"00",
													4283	=>X"00",
													4284	=>X"00",
													4285	=>X"00",
													4286	=>X"00",
													4287	=>X"00",
													4288	=>X"00",
													4289	=>X"00",
													4290	=>X"00",
													4291	=>X"00",
													4292	=>X"00",
													4293	=>X"00",
													4294	=>X"00",
													4295	=>X"00",
													4296	=>X"00",
													4297	=>X"00",
													4298	=>X"00",
													4299	=>X"00",
													4300	=>X"00",
													4301	=>X"00",
													4302	=>X"00",
													4303	=>X"00",
													4304	=>X"00",
													4305	=>X"00",
													4306	=>X"00",
													4307	=>X"00",
													4308	=>X"00",
													4309	=>X"1f",
													4310	=>X"83",
													4311	=>X"c0",
													4312	=>X"00",
													4313	=>X"00",
													4314	=>X"e0",
													4315	=>X"fc",
													4316	=>X"00",
													4317	=>X"00",
													4318	=>X"00",
													4319	=>X"00",
													4320	=>X"00",
													4321	=>X"00",
													4322	=>X"00",
													4323	=>X"00",
													4324	=>X"00",
													4325	=>X"00",
													4326	=>X"00",
													4327	=>X"00",
													4328	=>X"00",
													4329	=>X"00",
													4330	=>X"00",
													4331	=>X"00",
													4332	=>X"00",
													4333	=>X"00",
													4334	=>X"00",
													4335	=>X"00",
													4336	=>X"00",
													4337	=>X"00",
													4338	=>X"00",
													4339	=>X"00",
													4340	=>X"00",
													4341	=>X"00",
													4342	=>X"00",
													4343	=>X"00",
													4344	=>X"00",
													4345	=>X"00",
													4346	=>X"00",
													4347	=>X"00",
													4348	=>X"00",
													4349	=>X"1f",
													4350	=>X"83",
													4351	=>X"c0",
													4352	=>X"00",
													4353	=>X"00",
													4354	=>X"f0",
													4355	=>X"7c",
													4356	=>X"00",
													4357	=>X"00",
													4358	=>X"00",
													4359	=>X"00",
													4360	=>X"00",
													4361	=>X"00",
													4362	=>X"00",
													4363	=>X"00",
													4364	=>X"00",
													4365	=>X"00",
													4366	=>X"00",
													4367	=>X"00",
													4368	=>X"00",
													4369	=>X"00",
													4370	=>X"00",
													4371	=>X"00",
													4372	=>X"00",
													4373	=>X"00",
													4374	=>X"00",
													4375	=>X"00",
													4376	=>X"00",
													4377	=>X"00",
													4378	=>X"00",
													4379	=>X"00",
													4380	=>X"00",
													4381	=>X"00",
													4382	=>X"00",
													4383	=>X"00",
													4384	=>X"00",
													4385	=>X"00",
													4386	=>X"00",
													4387	=>X"00",
													4388	=>X"00",
													4389	=>X"1f",
													4390	=>X"83",
													4391	=>X"e0",
													4392	=>X"00",
													4393	=>X"00",
													4394	=>X"f0",
													4395	=>X"7c",
													4396	=>X"00",
													4397	=>X"00",
													4398	=>X"00",
													4399	=>X"00",
													4400	=>X"00",
													4401	=>X"00",
													4402	=>X"00",
													4403	=>X"00",
													4404	=>X"00",
													4405	=>X"00",
													4406	=>X"00",
													4407	=>X"00",
													4408	=>X"00",
													4409	=>X"00",
													4410	=>X"00",
													4411	=>X"00",
													4412	=>X"00",
													4413	=>X"00",
													4414	=>X"00",
													4415	=>X"00",
													4416	=>X"00",
													4417	=>X"00",
													4418	=>X"00",
													4419	=>X"00",
													4420	=>X"00",
													4421	=>X"00",
													4422	=>X"00",
													4423	=>X"00",
													4424	=>X"00",
													4425	=>X"00",
													4426	=>X"00",
													4427	=>X"00",
													4428	=>X"00",
													4429	=>X"1f",
													4430	=>X"83",
													4431	=>X"f0",
													4432	=>X"00",
													4433	=>X"00",
													4434	=>X"f0",
													4435	=>X"7c",
													4436	=>X"00",
													4437	=>X"00",
													4438	=>X"00",
													4439	=>X"00",
													4440	=>X"00",
													4441	=>X"00",
													4442	=>X"00",
													4443	=>X"00",
													4444	=>X"00",
													4445	=>X"00",
													4446	=>X"00",
													4447	=>X"00",
													4448	=>X"00",
													4449	=>X"00",
													4450	=>X"00",
													4451	=>X"00",
													4452	=>X"00",
													4453	=>X"00",
													4454	=>X"00",
													4455	=>X"00",
													4456	=>X"00",
													4457	=>X"00",
													4458	=>X"00",
													4459	=>X"00",
													4460	=>X"00",
													4461	=>X"00",
													4462	=>X"00",
													4463	=>X"00",
													4464	=>X"00",
													4465	=>X"00",
													4466	=>X"00",
													4467	=>X"00",
													4468	=>X"00",
													4469	=>X"1f",
													4470	=>X"03",
													4471	=>X"f8",
													4472	=>X"00",
													4473	=>X"01",
													4474	=>X"f0",
													4475	=>X"7c",
													4476	=>X"00",
													4477	=>X"00",
													4478	=>X"00",
													4479	=>X"00",
													4480	=>X"00",
													4481	=>X"00",
													4482	=>X"00",
													4483	=>X"00",
													4484	=>X"00",
													4485	=>X"00",
													4486	=>X"00",
													4487	=>X"00",
													4488	=>X"00",
													4489	=>X"00",
													4490	=>X"00",
													4491	=>X"00",
													4492	=>X"00",
													4493	=>X"00",
													4494	=>X"00",
													4495	=>X"00",
													4496	=>X"00",
													4497	=>X"00",
													4498	=>X"00",
													4499	=>X"00",
													4500	=>X"00",
													4501	=>X"00",
													4502	=>X"00",
													4503	=>X"00",
													4504	=>X"00",
													4505	=>X"00",
													4506	=>X"00",
													4507	=>X"00",
													4508	=>X"00",
													4509	=>X"1f",
													4510	=>X"00",
													4511	=>X"fc",
													4512	=>X"00",
													4513	=>X"03",
													4514	=>X"f0",
													4515	=>X"7c",
													4516	=>X"00",
													4517	=>X"00",
													4518	=>X"00",
													4519	=>X"00",
													4520	=>X"00",
													4521	=>X"00",
													4522	=>X"00",
													4523	=>X"00",
													4524	=>X"00",
													4525	=>X"00",
													4526	=>X"00",
													4527	=>X"00",
													4528	=>X"00",
													4529	=>X"00",
													4530	=>X"00",
													4531	=>X"00",
													4532	=>X"00",
													4533	=>X"00",
													4534	=>X"00",
													4535	=>X"00",
													4536	=>X"00",
													4537	=>X"00",
													4538	=>X"00",
													4539	=>X"00",
													4540	=>X"00",
													4541	=>X"00",
													4542	=>X"00",
													4543	=>X"00",
													4544	=>X"00",
													4545	=>X"00",
													4546	=>X"00",
													4547	=>X"00",
													4548	=>X"00",
													4549	=>X"1f",
													4550	=>X"00",
													4551	=>X"3f",
													4552	=>X"00",
													4553	=>X"0f",
													4554	=>X"f0",
													4555	=>X"7c",
													4556	=>X"00",
													4557	=>X"00",
													4558	=>X"00",
													4559	=>X"00",
													4560	=>X"00",
													4561	=>X"00",
													4562	=>X"00",
													4563	=>X"00",
													4564	=>X"00",
													4565	=>X"00",
													4566	=>X"00",
													4567	=>X"00",
													4568	=>X"00",
													4569	=>X"00",
													4570	=>X"00",
													4571	=>X"00",
													4572	=>X"00",
													4573	=>X"00",
													4574	=>X"00",
													4575	=>X"00",
													4576	=>X"00",
													4577	=>X"00",
													4578	=>X"00",
													4579	=>X"00",
													4580	=>X"00",
													4581	=>X"00",
													4582	=>X"00",
													4583	=>X"00",
													4584	=>X"00",
													4585	=>X"00",
													4586	=>X"00",
													4587	=>X"00",
													4588	=>X"00",
													4589	=>X"1f",
													4590	=>X"00",
													4591	=>X"0e",
													4592	=>X"00",
													4593	=>X"1f",
													4594	=>X"f0",
													4595	=>X"7c",
													4596	=>X"00",
													4597	=>X"00",
													4598	=>X"00",
													4599	=>X"00",
													4600	=>X"00",
													4601	=>X"00",
													4602	=>X"00",
													4603	=>X"00",
													4604	=>X"00",
													4605	=>X"00",
													4606	=>X"00",
													4607	=>X"00",
													4608	=>X"00",
													4609	=>X"00",
													4610	=>X"00",
													4611	=>X"00",
													4612	=>X"00",
													4613	=>X"00",
													4614	=>X"00",
													4615	=>X"00",
													4616	=>X"00",
													4617	=>X"00",
													4618	=>X"00",
													4619	=>X"00",
													4620	=>X"00",
													4621	=>X"00",
													4622	=>X"00",
													4623	=>X"00",
													4624	=>X"00",
													4625	=>X"00",
													4626	=>X"00",
													4627	=>X"00",
													4628	=>X"00",
													4629	=>X"1f",
													4630	=>X"03",
													4631	=>X"00",
													4632	=>X"00",
													4633	=>X"1f",
													4634	=>X"f0",
													4635	=>X"7c",
													4636	=>X"00",
													4637	=>X"00",
													4638	=>X"00",
													4639	=>X"00",
													4640	=>X"00",
													4641	=>X"00",
													4642	=>X"00",
													4643	=>X"00",
													4644	=>X"00",
													4645	=>X"00",
													4646	=>X"00",
													4647	=>X"00",
													4648	=>X"00",
													4649	=>X"00",
													4650	=>X"00",
													4651	=>X"00",
													4652	=>X"00",
													4653	=>X"00",
													4654	=>X"00",
													4655	=>X"00",
													4656	=>X"00",
													4657	=>X"00",
													4658	=>X"00",
													4659	=>X"00",
													4660	=>X"00",
													4661	=>X"00",
													4662	=>X"00",
													4663	=>X"00",
													4664	=>X"00",
													4665	=>X"00",
													4666	=>X"00",
													4667	=>X"00",
													4668	=>X"00",
													4669	=>X"1f",
													4670	=>X"03",
													4671	=>X"80",
													4672	=>X"00",
													4673	=>X"00",
													4674	=>X"00",
													4675	=>X"7c",
													4676	=>X"00",
													4677	=>X"00",
													4678	=>X"00",
													4679	=>X"00",
													4680	=>X"00",
													4681	=>X"00",
													4682	=>X"00",
													4683	=>X"00",
													4684	=>X"00",
													4685	=>X"00",
													4686	=>X"00",
													4687	=>X"00",
													4688	=>X"00",
													4689	=>X"00",
													4690	=>X"00",
													4691	=>X"00",
													4692	=>X"00",
													4693	=>X"00",
													4694	=>X"00",
													4695	=>X"00",
													4696	=>X"00",
													4697	=>X"00",
													4698	=>X"00",
													4699	=>X"00",
													4700	=>X"00",
													4701	=>X"00",
													4702	=>X"00",
													4703	=>X"00",
													4704	=>X"00",
													4705	=>X"00",
													4706	=>X"00",
													4707	=>X"00",
													4708	=>X"00",
													4709	=>X"1f",
													4710	=>X"03",
													4711	=>X"f0",
													4712	=>X"00",
													4713	=>X"00",
													4714	=>X"00",
													4715	=>X"7c",
													4716	=>X"00",
													4717	=>X"00",
													4718	=>X"00",
													4719	=>X"00",
													4720	=>X"00",
													4721	=>X"00",
													4722	=>X"00",
													4723	=>X"00",
													4724	=>X"00",
													4725	=>X"00",
													4726	=>X"00",
													4727	=>X"00",
													4728	=>X"00",
													4729	=>X"00",
													4730	=>X"00",
													4731	=>X"00",
													4732	=>X"00",
													4733	=>X"00",
													4734	=>X"00",
													4735	=>X"00",
													4736	=>X"00",
													4737	=>X"00",
													4738	=>X"00",
													4739	=>X"00",
													4740	=>X"00",
													4741	=>X"00",
													4742	=>X"00",
													4743	=>X"00",
													4744	=>X"00",
													4745	=>X"00",
													4746	=>X"00",
													4747	=>X"00",
													4748	=>X"00",
													4749	=>X"1f",
													4750	=>X"03",
													4751	=>X"ff",
													4752	=>X"00",
													4753	=>X"00",
													4754	=>X"00",
													4755	=>X"7c",
													4756	=>X"00",
													4757	=>X"00",
													4758	=>X"00",
													4759	=>X"00",
													4760	=>X"00",
													4761	=>X"00",
													4762	=>X"00",
													4763	=>X"00",
													4764	=>X"00",
													4765	=>X"00",
													4766	=>X"00",
													4767	=>X"00",
													4768	=>X"00",
													4769	=>X"00",
													4770	=>X"00",
													4771	=>X"00",
													4772	=>X"00",
													4773	=>X"00",
													4774	=>X"00",
													4775	=>X"00",
													4776	=>X"00",
													4777	=>X"00",
													4778	=>X"00",
													4779	=>X"00",
													4780	=>X"00",
													4781	=>X"00",
													4782	=>X"00",
													4783	=>X"00",
													4784	=>X"00",
													4785	=>X"00",
													4786	=>X"00",
													4787	=>X"00",
													4788	=>X"00",
													4789	=>X"1f",
													4790	=>X"03",
													4791	=>X"ff",
													4792	=>X"f0",
													4793	=>X"00",
													4794	=>X"00",
													4795	=>X"7c",
													4796	=>X"00",
													4797	=>X"00",
													4798	=>X"00",
													4799	=>X"00",
													4800	=>X"00",
													4801	=>X"00",
													4802	=>X"00",
													4803	=>X"00",
													4804	=>X"00",
													4805	=>X"00",
													4806	=>X"00",
													4807	=>X"00",
													4808	=>X"00",
													4809	=>X"00",
													4810	=>X"00",
													4811	=>X"00",
													4812	=>X"00",
													4813	=>X"00",
													4814	=>X"00",
													4815	=>X"00",
													4816	=>X"00",
													4817	=>X"00",
													4818	=>X"00",
													4819	=>X"00",
													4820	=>X"00",
													4821	=>X"00",
													4822	=>X"00",
													4823	=>X"00",
													4824	=>X"00",
													4825	=>X"00",
													4826	=>X"00",
													4827	=>X"00",
													4828	=>X"00",
													4829	=>X"1f",
													4830	=>X"03",
													4831	=>X"ff",
													4832	=>X"ff",
													4833	=>X"80",
													4834	=>X"00",
													4835	=>X"7c",
													4836	=>X"00",
													4837	=>X"00",
													4838	=>X"00",
													4839	=>X"00",
													4840	=>X"00",
													4841	=>X"00",
													4842	=>X"00",
													4843	=>X"00",
													4844	=>X"00",
													4845	=>X"00",
													4846	=>X"00",
													4847	=>X"00",
													4848	=>X"00",
													4849	=>X"00",
													4850	=>X"00",
													4851	=>X"00",
													4852	=>X"00",
													4853	=>X"00",
													4854	=>X"00",
													4855	=>X"00",
													4856	=>X"00",
													4857	=>X"00",
													4858	=>X"00",
													4859	=>X"00",
													4860	=>X"00",
													4861	=>X"00",
													4862	=>X"00",
													4863	=>X"00",
													4864	=>X"00",
													4865	=>X"00",
													4866	=>X"00",
													4867	=>X"00",
													4868	=>X"00",
													4869	=>X"1f",
													4870	=>X"03",
													4871	=>X"ff",
													4872	=>X"ff",
													4873	=>X"fc",
													4874	=>X"30",
													4875	=>X"7c",
													4876	=>X"00",
													4877	=>X"00",
													4878	=>X"00",
													4879	=>X"00",
													4880	=>X"00",
													4881	=>X"00",
													4882	=>X"00",
													4883	=>X"00",
													4884	=>X"00",
													4885	=>X"00",
													4886	=>X"00",
													4887	=>X"00",
													4888	=>X"00",
													4889	=>X"00",
													4890	=>X"00",
													4891	=>X"00",
													4892	=>X"00",
													4893	=>X"00",
													4894	=>X"00",
													4895	=>X"00",
													4896	=>X"00",
													4897	=>X"00",
													4898	=>X"00",
													4899	=>X"00",
													4900	=>X"00",
													4901	=>X"00",
													4902	=>X"00",
													4903	=>X"00",
													4904	=>X"00",
													4905	=>X"00",
													4906	=>X"00",
													4907	=>X"00",
													4908	=>X"00",
													4909	=>X"1f",
													4910	=>X"03",
													4911	=>X"8f",
													4912	=>X"ff",
													4913	=>X"ff",
													4914	=>X"f0",
													4915	=>X"fc",
													4916	=>X"00",
													4917	=>X"00",
													4918	=>X"00",
													4919	=>X"00",
													4920	=>X"00",
													4921	=>X"00",
													4922	=>X"00",
													4923	=>X"00",
													4924	=>X"00",
													4925	=>X"00",
													4926	=>X"00",
													4927	=>X"00",
													4928	=>X"00",
													4929	=>X"00",
													4930	=>X"00",
													4931	=>X"00",
													4932	=>X"00",
													4933	=>X"00",
													4934	=>X"00",
													4935	=>X"00",
													4936	=>X"00",
													4937	=>X"00",
													4938	=>X"00",
													4939	=>X"00",
													4940	=>X"00",
													4941	=>X"00",
													4942	=>X"00",
													4943	=>X"00",
													4944	=>X"00",
													4945	=>X"00",
													4946	=>X"00",
													4947	=>X"00",
													4948	=>X"00",
													4949	=>X"1f",
													4950	=>X"00",
													4951	=>X"00",
													4952	=>X"ff",
													4953	=>X"ff",
													4954	=>X"f0",
													4955	=>X"fc",
													4956	=>X"00",
													4957	=>X"00",
													4958	=>X"00",
													4959	=>X"00",
													4960	=>X"00",
													4961	=>X"00",
													4962	=>X"00",
													4963	=>X"00",
													4964	=>X"00",
													4965	=>X"00",
													4966	=>X"00",
													4967	=>X"00",
													4968	=>X"00",
													4969	=>X"00",
													4970	=>X"00",
													4971	=>X"00",
													4972	=>X"00",
													4973	=>X"00",
													4974	=>X"00",
													4975	=>X"00",
													4976	=>X"00",
													4977	=>X"00",
													4978	=>X"00",
													4979	=>X"00",
													4980	=>X"00",
													4981	=>X"00",
													4982	=>X"00",
													4983	=>X"00",
													4984	=>X"00",
													4985	=>X"00",
													4986	=>X"00",
													4987	=>X"00",
													4988	=>X"00",
													4989	=>X"1f",
													4990	=>X"00",
													4991	=>X"00",
													4992	=>X"3f",
													4993	=>X"ff",
													4994	=>X"f0",
													4995	=>X"fc",
													4996	=>X"00",
													4997	=>X"00",
													4998	=>X"00",
													4999	=>X"00",
													5000	=>X"00",
													5001	=>X"00",
													5002	=>X"00",
													5003	=>X"00",
													5004	=>X"00",
													5005	=>X"00",
													5006	=>X"00",
													5007	=>X"00",
													5008	=>X"00",
													5009	=>X"00",
													5010	=>X"00",
													5011	=>X"00",
													5012	=>X"00",
													5013	=>X"00",
													5014	=>X"00",
													5015	=>X"00",
													5016	=>X"00",
													5017	=>X"00",
													5018	=>X"00",
													5019	=>X"00",
													5020	=>X"00",
													5021	=>X"00",
													5022	=>X"00",
													5023	=>X"00",
													5024	=>X"00",
													5025	=>X"00",
													5026	=>X"00",
													5027	=>X"00",
													5028	=>X"00",
													5029	=>X"1f",
													5030	=>X"80",
													5031	=>X"00",
													5032	=>X"1e",
													5033	=>X"7f",
													5034	=>X"f0",
													5035	=>X"fc",
													5036	=>X"00",
													5037	=>X"00",
													5038	=>X"00",
													5039	=>X"00",
													5040	=>X"00",
													5041	=>X"00",
													5042	=>X"00",
													5043	=>X"00",
													5044	=>X"00",
													5045	=>X"00",
													5046	=>X"00",
													5047	=>X"00",
													5048	=>X"00",
													5049	=>X"00",
													5050	=>X"00",
													5051	=>X"00",
													5052	=>X"00",
													5053	=>X"00",
													5054	=>X"00",
													5055	=>X"00",
													5056	=>X"00",
													5057	=>X"00",
													5058	=>X"00",
													5059	=>X"00",
													5060	=>X"00",
													5061	=>X"00",
													5062	=>X"00",
													5063	=>X"00",
													5064	=>X"00",
													5065	=>X"00",
													5066	=>X"00",
													5067	=>X"00",
													5068	=>X"00",
													5069	=>X"1f",
													5070	=>X"80",
													5071	=>X"00",
													5072	=>X"0f",
													5073	=>X"03",
													5074	=>X"f0",
													5075	=>X"fc",
													5076	=>X"00",
													5077	=>X"00",
													5078	=>X"00",
													5079	=>X"00",
													5080	=>X"00",
													5081	=>X"00",
													5082	=>X"00",
													5083	=>X"00",
													5084	=>X"00",
													5085	=>X"00",
													5086	=>X"00",
													5087	=>X"00",
													5088	=>X"00",
													5089	=>X"00",
													5090	=>X"00",
													5091	=>X"00",
													5092	=>X"00",
													5093	=>X"00",
													5094	=>X"00",
													5095	=>X"00",
													5096	=>X"00",
													5097	=>X"00",
													5098	=>X"00",
													5099	=>X"00",
													5100	=>X"00",
													5101	=>X"00",
													5102	=>X"00",
													5103	=>X"00",
													5104	=>X"00",
													5105	=>X"00",
													5106	=>X"00",
													5107	=>X"00",
													5108	=>X"00",
													5109	=>X"1f",
													5110	=>X"80",
													5111	=>X"00",
													5112	=>X"07",
													5113	=>X"80",
													5114	=>X"f0",
													5115	=>X"fc",
													5116	=>X"00",
													5117	=>X"00",
													5118	=>X"00",
													5119	=>X"00",
													5120	=>X"00",
													5121	=>X"00",
													5122	=>X"00",
													5123	=>X"00",
													5124	=>X"00",
													5125	=>X"00",
													5126	=>X"00",
													5127	=>X"00",
													5128	=>X"00",
													5129	=>X"00",
													5130	=>X"00",
													5131	=>X"00",
													5132	=>X"00",
													5133	=>X"00",
													5134	=>X"00",
													5135	=>X"00",
													5136	=>X"00",
													5137	=>X"00",
													5138	=>X"00",
													5139	=>X"00",
													5140	=>X"00",
													5141	=>X"00",
													5142	=>X"00",
													5143	=>X"00",
													5144	=>X"00",
													5145	=>X"00",
													5146	=>X"00",
													5147	=>X"00",
													5148	=>X"00",
													5149	=>X"1f",
													5150	=>X"83",
													5151	=>X"00",
													5152	=>X"03",
													5153	=>X"c0",
													5154	=>X"30",
													5155	=>X"fc",
													5156	=>X"00",
													5157	=>X"00",
													5158	=>X"00",
													5159	=>X"00",
													5160	=>X"00",
													5161	=>X"00",
													5162	=>X"00",
													5163	=>X"00",
													5164	=>X"00",
													5165	=>X"00",
													5166	=>X"00",
													5167	=>X"00",
													5168	=>X"00",
													5169	=>X"00",
													5170	=>X"00",
													5171	=>X"00",
													5172	=>X"00",
													5173	=>X"00",
													5174	=>X"00",
													5175	=>X"00",
													5176	=>X"00",
													5177	=>X"00",
													5178	=>X"00",
													5179	=>X"00",
													5180	=>X"00",
													5181	=>X"00",
													5182	=>X"00",
													5183	=>X"00",
													5184	=>X"00",
													5185	=>X"00",
													5186	=>X"00",
													5187	=>X"00",
													5188	=>X"00",
													5189	=>X"1f",
													5190	=>X"83",
													5191	=>X"80",
													5192	=>X"01",
													5193	=>X"e0",
													5194	=>X"20",
													5195	=>X"fc",
													5196	=>X"00",
													5197	=>X"00",
													5198	=>X"00",
													5199	=>X"00",
													5200	=>X"00",
													5201	=>X"00",
													5202	=>X"00",
													5203	=>X"00",
													5204	=>X"00",
													5205	=>X"00",
													5206	=>X"00",
													5207	=>X"00",
													5208	=>X"00",
													5209	=>X"00",
													5210	=>X"00",
													5211	=>X"00",
													5212	=>X"00",
													5213	=>X"00",
													5214	=>X"00",
													5215	=>X"00",
													5216	=>X"00",
													5217	=>X"00",
													5218	=>X"00",
													5219	=>X"00",
													5220	=>X"00",
													5221	=>X"00",
													5222	=>X"00",
													5223	=>X"00",
													5224	=>X"00",
													5225	=>X"00",
													5226	=>X"00",
													5227	=>X"00",
													5228	=>X"00",
													5229	=>X"1f",
													5230	=>X"83",
													5231	=>X"f0",
													5232	=>X"01",
													5233	=>X"f0",
													5234	=>X"00",
													5235	=>X"fc",
													5236	=>X"00",
													5237	=>X"00",
													5238	=>X"00",
													5239	=>X"00",
													5240	=>X"00",
													5241	=>X"00",
													5242	=>X"00",
													5243	=>X"00",
													5244	=>X"00",
													5245	=>X"00",
													5246	=>X"00",
													5247	=>X"00",
													5248	=>X"00",
													5249	=>X"00",
													5250	=>X"00",
													5251	=>X"00",
													5252	=>X"00",
													5253	=>X"00",
													5254	=>X"00",
													5255	=>X"00",
													5256	=>X"00",
													5257	=>X"00",
													5258	=>X"00",
													5259	=>X"00",
													5260	=>X"00",
													5261	=>X"00",
													5262	=>X"00",
													5263	=>X"00",
													5264	=>X"00",
													5265	=>X"00",
													5266	=>X"00",
													5267	=>X"00",
													5268	=>X"00",
													5269	=>X"1f",
													5270	=>X"83",
													5271	=>X"ff",
													5272	=>X"00",
													5273	=>X"f8",
													5274	=>X"00",
													5275	=>X"f8",
													5276	=>X"00",
													5277	=>X"00",
													5278	=>X"00",
													5279	=>X"00",
													5280	=>X"00",
													5281	=>X"00",
													5282	=>X"00",
													5283	=>X"00",
													5284	=>X"00",
													5285	=>X"00",
													5286	=>X"00",
													5287	=>X"00",
													5288	=>X"00",
													5289	=>X"00",
													5290	=>X"00",
													5291	=>X"00",
													5292	=>X"00",
													5293	=>X"00",
													5294	=>X"00",
													5295	=>X"00",
													5296	=>X"00",
													5297	=>X"00",
													5298	=>X"00",
													5299	=>X"00",
													5300	=>X"00",
													5301	=>X"00",
													5302	=>X"00",
													5303	=>X"00",
													5304	=>X"00",
													5305	=>X"00",
													5306	=>X"00",
													5307	=>X"00",
													5308	=>X"00",
													5309	=>X"1f",
													5310	=>X"83",
													5311	=>X"ff",
													5312	=>X"f0",
													5313	=>X"7c",
													5314	=>X"00",
													5315	=>X"f8",
													5316	=>X"00",
													5317	=>X"00",
													5318	=>X"00",
													5319	=>X"00",
													5320	=>X"00",
													5321	=>X"00",
													5322	=>X"00",
													5323	=>X"00",
													5324	=>X"00",
													5325	=>X"00",
													5326	=>X"00",
													5327	=>X"00",
													5328	=>X"00",
													5329	=>X"00",
													5330	=>X"00",
													5331	=>X"00",
													5332	=>X"00",
													5333	=>X"00",
													5334	=>X"00",
													5335	=>X"00",
													5336	=>X"00",
													5337	=>X"00",
													5338	=>X"00",
													5339	=>X"00",
													5340	=>X"00",
													5341	=>X"00",
													5342	=>X"00",
													5343	=>X"00",
													5344	=>X"00",
													5345	=>X"00",
													5346	=>X"00",
													5347	=>X"00",
													5348	=>X"00",
													5349	=>X"0f",
													5350	=>X"83",
													5351	=>X"ff",
													5352	=>X"ff",
													5353	=>X"bc",
													5354	=>X"00",
													5355	=>X"f8",
													5356	=>X"00",
													5357	=>X"00",
													5358	=>X"00",
													5359	=>X"00",
													5360	=>X"00",
													5361	=>X"00",
													5362	=>X"00",
													5363	=>X"00",
													5364	=>X"00",
													5365	=>X"00",
													5366	=>X"00",
													5367	=>X"00",
													5368	=>X"00",
													5369	=>X"00",
													5370	=>X"00",
													5371	=>X"00",
													5372	=>X"00",
													5373	=>X"00",
													5374	=>X"00",
													5375	=>X"00",
													5376	=>X"00",
													5377	=>X"00",
													5378	=>X"00",
													5379	=>X"00",
													5380	=>X"00",
													5381	=>X"00",
													5382	=>X"00",
													5383	=>X"00",
													5384	=>X"00",
													5385	=>X"00",
													5386	=>X"00",
													5387	=>X"00",
													5388	=>X"00",
													5389	=>X"0f",
													5390	=>X"83",
													5391	=>X"ff",
													5392	=>X"ff",
													5393	=>X"fe",
													5394	=>X"70",
													5395	=>X"f8",
													5396	=>X"00",
													5397	=>X"00",
													5398	=>X"00",
													5399	=>X"00",
													5400	=>X"00",
													5401	=>X"00",
													5402	=>X"00",
													5403	=>X"00",
													5404	=>X"00",
													5405	=>X"00",
													5406	=>X"00",
													5407	=>X"00",
													5408	=>X"00",
													5409	=>X"00",
													5410	=>X"00",
													5411	=>X"00",
													5412	=>X"00",
													5413	=>X"00",
													5414	=>X"00",
													5415	=>X"00",
													5416	=>X"00",
													5417	=>X"00",
													5418	=>X"00",
													5419	=>X"00",
													5420	=>X"00",
													5421	=>X"00",
													5422	=>X"00",
													5423	=>X"00",
													5424	=>X"00",
													5425	=>X"00",
													5426	=>X"00",
													5427	=>X"00",
													5428	=>X"00",
													5429	=>X"0f",
													5430	=>X"83",
													5431	=>X"8f",
													5432	=>X"ff",
													5433	=>X"ff",
													5434	=>X"f0",
													5435	=>X"f8",
													5436	=>X"00",
													5437	=>X"00",
													5438	=>X"00",
													5439	=>X"00",
													5440	=>X"00",
													5441	=>X"00",
													5442	=>X"00",
													5443	=>X"00",
													5444	=>X"00",
													5445	=>X"00",
													5446	=>X"00",
													5447	=>X"00",
													5448	=>X"00",
													5449	=>X"00",
													5450	=>X"00",
													5451	=>X"00",
													5452	=>X"00",
													5453	=>X"00",
													5454	=>X"00",
													5455	=>X"00",
													5456	=>X"00",
													5457	=>X"00",
													5458	=>X"00",
													5459	=>X"00",
													5460	=>X"00",
													5461	=>X"00",
													5462	=>X"00",
													5463	=>X"00",
													5464	=>X"00",
													5465	=>X"00",
													5466	=>X"00",
													5467	=>X"00",
													5468	=>X"00",
													5469	=>X"0f",
													5470	=>X"81",
													5471	=>X"00",
													5472	=>X"7f",
													5473	=>X"ff",
													5474	=>X"f0",
													5475	=>X"f8",
													5476	=>X"00",
													5477	=>X"00",
													5478	=>X"00",
													5479	=>X"00",
													5480	=>X"00",
													5481	=>X"00",
													5482	=>X"00",
													5483	=>X"00",
													5484	=>X"00",
													5485	=>X"00",
													5486	=>X"00",
													5487	=>X"00",
													5488	=>X"00",
													5489	=>X"00",
													5490	=>X"00",
													5491	=>X"00",
													5492	=>X"00",
													5493	=>X"00",
													5494	=>X"00",
													5495	=>X"00",
													5496	=>X"00",
													5497	=>X"00",
													5498	=>X"00",
													5499	=>X"00",
													5500	=>X"00",
													5501	=>X"00",
													5502	=>X"00",
													5503	=>X"00",
													5504	=>X"00",
													5505	=>X"00",
													5506	=>X"00",
													5507	=>X"00",
													5508	=>X"00",
													5509	=>X"0f",
													5510	=>X"80",
													5511	=>X"00",
													5512	=>X"07",
													5513	=>X"ff",
													5514	=>X"f0",
													5515	=>X"f8",
													5516	=>X"00",
													5517	=>X"00",
													5518	=>X"00",
													5519	=>X"00",
													5520	=>X"00",
													5521	=>X"00",
													5522	=>X"00",
													5523	=>X"00",
													5524	=>X"00",
													5525	=>X"00",
													5526	=>X"00",
													5527	=>X"00",
													5528	=>X"00",
													5529	=>X"00",
													5530	=>X"00",
													5531	=>X"00",
													5532	=>X"00",
													5533	=>X"00",
													5534	=>X"00",
													5535	=>X"00",
													5536	=>X"00",
													5537	=>X"00",
													5538	=>X"00",
													5539	=>X"00",
													5540	=>X"00",
													5541	=>X"00",
													5542	=>X"00",
													5543	=>X"00",
													5544	=>X"00",
													5545	=>X"00",
													5546	=>X"00",
													5547	=>X"00",
													5548	=>X"00",
													5549	=>X"0f",
													5550	=>X"80",
													5551	=>X"00",
													5552	=>X"00",
													5553	=>X"7f",
													5554	=>X"f0",
													5555	=>X"f8",
													5556	=>X"00",
													5557	=>X"00",
													5558	=>X"00",
													5559	=>X"00",
													5560	=>X"00",
													5561	=>X"00",
													5562	=>X"00",
													5563	=>X"00",
													5564	=>X"00",
													5565	=>X"00",
													5566	=>X"00",
													5567	=>X"00",
													5568	=>X"00",
													5569	=>X"00",
													5570	=>X"00",
													5571	=>X"00",
													5572	=>X"00",
													5573	=>X"00",
													5574	=>X"00",
													5575	=>X"00",
													5576	=>X"00",
													5577	=>X"00",
													5578	=>X"00",
													5579	=>X"00",
													5580	=>X"00",
													5581	=>X"00",
													5582	=>X"00",
													5583	=>X"00",
													5584	=>X"00",
													5585	=>X"00",
													5586	=>X"00",
													5587	=>X"00",
													5588	=>X"00",
													5589	=>X"0f",
													5590	=>X"80",
													5591	=>X"00",
													5592	=>X"00",
													5593	=>X"07",
													5594	=>X"f0",
													5595	=>X"f8",
													5596	=>X"00",
													5597	=>X"00",
													5598	=>X"00",
													5599	=>X"00",
													5600	=>X"00",
													5601	=>X"00",
													5602	=>X"00",
													5603	=>X"00",
													5604	=>X"00",
													5605	=>X"00",
													5606	=>X"00",
													5607	=>X"00",
													5608	=>X"00",
													5609	=>X"00",
													5610	=>X"00",
													5611	=>X"00",
													5612	=>X"00",
													5613	=>X"00",
													5614	=>X"00",
													5615	=>X"00",
													5616	=>X"00",
													5617	=>X"00",
													5618	=>X"00",
													5619	=>X"00",
													5620	=>X"00",
													5621	=>X"00",
													5622	=>X"00",
													5623	=>X"00",
													5624	=>X"00",
													5625	=>X"00",
													5626	=>X"00",
													5627	=>X"00",
													5628	=>X"00",
													5629	=>X"0f",
													5630	=>X"83",
													5631	=>X"ff",
													5632	=>X"00",
													5633	=>X"00",
													5634	=>X"f1",
													5635	=>X"f8",
													5636	=>X"00",
													5637	=>X"00",
													5638	=>X"00",
													5639	=>X"00",
													5640	=>X"00",
													5641	=>X"00",
													5642	=>X"00",
													5643	=>X"00",
													5644	=>X"00",
													5645	=>X"00",
													5646	=>X"00",
													5647	=>X"00",
													5648	=>X"00",
													5649	=>X"00",
													5650	=>X"00",
													5651	=>X"00",
													5652	=>X"00",
													5653	=>X"00",
													5654	=>X"00",
													5655	=>X"00",
													5656	=>X"00",
													5657	=>X"00",
													5658	=>X"00",
													5659	=>X"00",
													5660	=>X"00",
													5661	=>X"00",
													5662	=>X"00",
													5663	=>X"00",
													5664	=>X"00",
													5665	=>X"00",
													5666	=>X"00",
													5667	=>X"00",
													5668	=>X"00",
													5669	=>X"0f",
													5670	=>X"83",
													5671	=>X"fc",
													5672	=>X"00",
													5673	=>X"00",
													5674	=>X"61",
													5675	=>X"f0",
													5676	=>X"00",
													5677	=>X"00",
													5678	=>X"00",
													5679	=>X"00",
													5680	=>X"00",
													5681	=>X"00",
													5682	=>X"00",
													5683	=>X"00",
													5684	=>X"00",
													5685	=>X"00",
													5686	=>X"00",
													5687	=>X"00",
													5688	=>X"00",
													5689	=>X"00",
													5690	=>X"00",
													5691	=>X"00",
													5692	=>X"00",
													5693	=>X"00",
													5694	=>X"00",
													5695	=>X"00",
													5696	=>X"00",
													5697	=>X"00",
													5698	=>X"00",
													5699	=>X"00",
													5700	=>X"00",
													5701	=>X"00",
													5702	=>X"00",
													5703	=>X"00",
													5704	=>X"00",
													5705	=>X"00",
													5706	=>X"00",
													5707	=>X"00",
													5708	=>X"00",
													5709	=>X"0f",
													5710	=>X"83",
													5711	=>X"f8",
													5712	=>X"00",
													5713	=>X"00",
													5714	=>X"21",
													5715	=>X"f0",
													5716	=>X"00",
													5717	=>X"00",
													5718	=>X"00",
													5719	=>X"00",
													5720	=>X"00",
													5721	=>X"00",
													5722	=>X"00",
													5723	=>X"00",
													5724	=>X"00",
													5725	=>X"00",
													5726	=>X"00",
													5727	=>X"00",
													5728	=>X"00",
													5729	=>X"00",
													5730	=>X"00",
													5731	=>X"00",
													5732	=>X"00",
													5733	=>X"00",
													5734	=>X"00",
													5735	=>X"00",
													5736	=>X"00",
													5737	=>X"00",
													5738	=>X"00",
													5739	=>X"00",
													5740	=>X"00",
													5741	=>X"00",
													5742	=>X"00",
													5743	=>X"00",
													5744	=>X"00",
													5745	=>X"00",
													5746	=>X"00",
													5747	=>X"00",
													5748	=>X"00",
													5749	=>X"0f",
													5750	=>X"81",
													5751	=>X"f0",
													5752	=>X"00",
													5753	=>X"00",
													5754	=>X"01",
													5755	=>X"f0",
													5756	=>X"00",
													5757	=>X"00",
													5758	=>X"00",
													5759	=>X"00",
													5760	=>X"00",
													5761	=>X"00",
													5762	=>X"00",
													5763	=>X"00",
													5764	=>X"00",
													5765	=>X"00",
													5766	=>X"00",
													5767	=>X"00",
													5768	=>X"00",
													5769	=>X"00",
													5770	=>X"00",
													5771	=>X"00",
													5772	=>X"00",
													5773	=>X"00",
													5774	=>X"00",
													5775	=>X"00",
													5776	=>X"00",
													5777	=>X"00",
													5778	=>X"00",
													5779	=>X"00",
													5780	=>X"00",
													5781	=>X"00",
													5782	=>X"00",
													5783	=>X"00",
													5784	=>X"00",
													5785	=>X"00",
													5786	=>X"00",
													5787	=>X"00",
													5788	=>X"00",
													5789	=>X"0f",
													5790	=>X"c1",
													5791	=>X"e0",
													5792	=>X"00",
													5793	=>X"1c",
													5794	=>X"01",
													5795	=>X"f0",
													5796	=>X"00",
													5797	=>X"00",
													5798	=>X"00",
													5799	=>X"00",
													5800	=>X"00",
													5801	=>X"00",
													5802	=>X"00",
													5803	=>X"00",
													5804	=>X"00",
													5805	=>X"00",
													5806	=>X"00",
													5807	=>X"00",
													5808	=>X"00",
													5809	=>X"00",
													5810	=>X"00",
													5811	=>X"00",
													5812	=>X"00",
													5813	=>X"00",
													5814	=>X"00",
													5815	=>X"00",
													5816	=>X"00",
													5817	=>X"00",
													5818	=>X"00",
													5819	=>X"00",
													5820	=>X"00",
													5821	=>X"00",
													5822	=>X"00",
													5823	=>X"00",
													5824	=>X"00",
													5825	=>X"00",
													5826	=>X"00",
													5827	=>X"00",
													5828	=>X"00",
													5829	=>X"0f",
													5830	=>X"c1",
													5831	=>X"e0",
													5832	=>X"00",
													5833	=>X"1e",
													5834	=>X"01",
													5835	=>X"f0",
													5836	=>X"00",
													5837	=>X"00",
													5838	=>X"00",
													5839	=>X"00",
													5840	=>X"00",
													5841	=>X"00",
													5842	=>X"00",
													5843	=>X"00",
													5844	=>X"00",
													5845	=>X"00",
													5846	=>X"00",
													5847	=>X"00",
													5848	=>X"00",
													5849	=>X"00",
													5850	=>X"00",
													5851	=>X"00",
													5852	=>X"00",
													5853	=>X"00",
													5854	=>X"00",
													5855	=>X"00",
													5856	=>X"00",
													5857	=>X"00",
													5858	=>X"00",
													5859	=>X"00",
													5860	=>X"00",
													5861	=>X"00",
													5862	=>X"00",
													5863	=>X"00",
													5864	=>X"00",
													5865	=>X"00",
													5866	=>X"00",
													5867	=>X"00",
													5868	=>X"00",
													5869	=>X"07",
													5870	=>X"c1",
													5871	=>X"c0",
													5872	=>X"00",
													5873	=>X"0f",
													5874	=>X"c1",
													5875	=>X"f0",
													5876	=>X"00",
													5877	=>X"00",
													5878	=>X"00",
													5879	=>X"00",
													5880	=>X"00",
													5881	=>X"00",
													5882	=>X"00",
													5883	=>X"00",
													5884	=>X"00",
													5885	=>X"00",
													5886	=>X"00",
													5887	=>X"00",
													5888	=>X"00",
													5889	=>X"00",
													5890	=>X"00",
													5891	=>X"00",
													5892	=>X"00",
													5893	=>X"00",
													5894	=>X"00",
													5895	=>X"00",
													5896	=>X"00",
													5897	=>X"00",
													5898	=>X"00",
													5899	=>X"00",
													5900	=>X"00",
													5901	=>X"00",
													5902	=>X"00",
													5903	=>X"00",
													5904	=>X"00",
													5905	=>X"00",
													5906	=>X"00",
													5907	=>X"00",
													5908	=>X"00",
													5909	=>X"07",
													5910	=>X"c1",
													5911	=>X"c0",
													5912	=>X"0f",
													5913	=>X"07",
													5914	=>X"e1",
													5915	=>X"f0",
													5916	=>X"00",
													5917	=>X"00",
													5918	=>X"00",
													5919	=>X"00",
													5920	=>X"00",
													5921	=>X"00",
													5922	=>X"00",
													5923	=>X"00",
													5924	=>X"00",
													5925	=>X"00",
													5926	=>X"00",
													5927	=>X"00",
													5928	=>X"00",
													5929	=>X"00",
													5930	=>X"00",
													5931	=>X"00",
													5932	=>X"00",
													5933	=>X"00",
													5934	=>X"00",
													5935	=>X"00",
													5936	=>X"00",
													5937	=>X"00",
													5938	=>X"00",
													5939	=>X"00",
													5940	=>X"00",
													5941	=>X"00",
													5942	=>X"00",
													5943	=>X"00",
													5944	=>X"00",
													5945	=>X"00",
													5946	=>X"00",
													5947	=>X"00",
													5948	=>X"00",
													5949	=>X"07",
													5950	=>X"c1",
													5951	=>X"e0",
													5952	=>X"0f",
													5953	=>X"03",
													5954	=>X"e3",
													5955	=>X"f0",
													5956	=>X"00",
													5957	=>X"00",
													5958	=>X"00",
													5959	=>X"00",
													5960	=>X"00",
													5961	=>X"00",
													5962	=>X"00",
													5963	=>X"00",
													5964	=>X"00",
													5965	=>X"00",
													5966	=>X"00",
													5967	=>X"00",
													5968	=>X"00",
													5969	=>X"00",
													5970	=>X"00",
													5971	=>X"00",
													5972	=>X"00",
													5973	=>X"00",
													5974	=>X"00",
													5975	=>X"00",
													5976	=>X"00",
													5977	=>X"00",
													5978	=>X"00",
													5979	=>X"00",
													5980	=>X"00",
													5981	=>X"00",
													5982	=>X"00",
													5983	=>X"00",
													5984	=>X"00",
													5985	=>X"00",
													5986	=>X"00",
													5987	=>X"00",
													5988	=>X"00",
													5989	=>X"07",
													5990	=>X"c1",
													5991	=>X"e0",
													5992	=>X"0f",
													5993	=>X"03",
													5994	=>X"e3",
													5995	=>X"f0",
													5996	=>X"00",
													5997	=>X"00",
													5998	=>X"00",
													5999	=>X"00",
													6000	=>X"00",
													6001	=>X"00",
													6002	=>X"00",
													6003	=>X"00",
													6004	=>X"00",
													6005	=>X"00",
													6006	=>X"00",
													6007	=>X"00",
													6008	=>X"00",
													6009	=>X"00",
													6010	=>X"00",
													6011	=>X"00",
													6012	=>X"00",
													6013	=>X"00",
													6014	=>X"00",
													6015	=>X"00",
													6016	=>X"00",
													6017	=>X"00",
													6018	=>X"00",
													6019	=>X"00",
													6020	=>X"00",
													6021	=>X"00",
													6022	=>X"00",
													6023	=>X"00",
													6024	=>X"00",
													6025	=>X"00",
													6026	=>X"00",
													6027	=>X"00",
													6028	=>X"00",
													6029	=>X"07",
													6030	=>X"c0",
													6031	=>X"f0",
													6032	=>X"0f",
													6033	=>X"01",
													6034	=>X"e3",
													6035	=>X"f0",
													6036	=>X"00",
													6037	=>X"00",
													6038	=>X"00",
													6039	=>X"00",
													6040	=>X"00",
													6041	=>X"00",
													6042	=>X"00",
													6043	=>X"00",
													6044	=>X"00",
													6045	=>X"00",
													6046	=>X"00",
													6047	=>X"00",
													6048	=>X"00",
													6049	=>X"00",
													6050	=>X"00",
													6051	=>X"00",
													6052	=>X"00",
													6053	=>X"00",
													6054	=>X"00",
													6055	=>X"00",
													6056	=>X"00",
													6057	=>X"00",
													6058	=>X"00",
													6059	=>X"00",
													6060	=>X"00",
													6061	=>X"00",
													6062	=>X"00",
													6063	=>X"00",
													6064	=>X"00",
													6065	=>X"00",
													6066	=>X"00",
													6067	=>X"00",
													6068	=>X"00",
													6069	=>X"07",
													6070	=>X"e0",
													6071	=>X"f8",
													6072	=>X"0f",
													6073	=>X"01",
													6074	=>X"c3",
													6075	=>X"e0",
													6076	=>X"00",
													6077	=>X"00",
													6078	=>X"00",
													6079	=>X"00",
													6080	=>X"00",
													6081	=>X"00",
													6082	=>X"00",
													6083	=>X"00",
													6084	=>X"00",
													6085	=>X"00",
													6086	=>X"00",
													6087	=>X"00",
													6088	=>X"00",
													6089	=>X"00",
													6090	=>X"00",
													6091	=>X"00",
													6092	=>X"00",
													6093	=>X"00",
													6094	=>X"00",
													6095	=>X"00",
													6096	=>X"00",
													6097	=>X"00",
													6098	=>X"00",
													6099	=>X"00",
													6100	=>X"00",
													6101	=>X"00",
													6102	=>X"00",
													6103	=>X"00",
													6104	=>X"00",
													6105	=>X"00",
													6106	=>X"00",
													6107	=>X"00",
													6108	=>X"00",
													6109	=>X"07",
													6110	=>X"e0",
													6111	=>X"f8",
													6112	=>X"0f",
													6113	=>X"01",
													6114	=>X"c3",
													6115	=>X"e0",
													6116	=>X"00",
													6117	=>X"00",
													6118	=>X"00",
													6119	=>X"00",
													6120	=>X"00",
													6121	=>X"00",
													6122	=>X"00",
													6123	=>X"00",
													6124	=>X"00",
													6125	=>X"00",
													6126	=>X"00",
													6127	=>X"00",
													6128	=>X"00",
													6129	=>X"00",
													6130	=>X"00",
													6131	=>X"00",
													6132	=>X"00",
													6133	=>X"00",
													6134	=>X"00",
													6135	=>X"00",
													6136	=>X"00",
													6137	=>X"00",
													6138	=>X"00",
													6139	=>X"00",
													6140	=>X"00",
													6141	=>X"00",
													6142	=>X"00",
													6143	=>X"00",
													6144	=>X"00",
													6145	=>X"00",
													6146	=>X"00",
													6147	=>X"00",
													6148	=>X"00",
													6149	=>X"07",
													6150	=>X"e0",
													6151	=>X"7c",
													6152	=>X"0f",
													6153	=>X"03",
													6154	=>X"c7",
													6155	=>X"e0",
													6156	=>X"00",
													6157	=>X"00",
													6158	=>X"00",
													6159	=>X"00",
													6160	=>X"00",
													6161	=>X"00",
													6162	=>X"00",
													6163	=>X"00",
													6164	=>X"00",
													6165	=>X"00",
													6166	=>X"00",
													6167	=>X"00",
													6168	=>X"00",
													6169	=>X"00",
													6170	=>X"00",
													6171	=>X"00",
													6172	=>X"00",
													6173	=>X"00",
													6174	=>X"00",
													6175	=>X"00",
													6176	=>X"00",
													6177	=>X"00",
													6178	=>X"00",
													6179	=>X"00",
													6180	=>X"00",
													6181	=>X"00",
													6182	=>X"00",
													6183	=>X"00",
													6184	=>X"00",
													6185	=>X"00",
													6186	=>X"00",
													6187	=>X"00",
													6188	=>X"00",
													6189	=>X"03",
													6190	=>X"e0",
													6191	=>X"7f",
													6192	=>X"0f",
													6193	=>X"07",
													6194	=>X"c7",
													6195	=>X"e0",
													6196	=>X"00",
													6197	=>X"00",
													6198	=>X"00",
													6199	=>X"00",
													6200	=>X"00",
													6201	=>X"00",
													6202	=>X"00",
													6203	=>X"00",
													6204	=>X"00",
													6205	=>X"00",
													6206	=>X"00",
													6207	=>X"00",
													6208	=>X"00",
													6209	=>X"00",
													6210	=>X"00",
													6211	=>X"00",
													6212	=>X"00",
													6213	=>X"00",
													6214	=>X"00",
													6215	=>X"00",
													6216	=>X"00",
													6217	=>X"00",
													6218	=>X"00",
													6219	=>X"00",
													6220	=>X"00",
													6221	=>X"00",
													6222	=>X"00",
													6223	=>X"00",
													6224	=>X"00",
													6225	=>X"00",
													6226	=>X"00",
													6227	=>X"00",
													6228	=>X"00",
													6229	=>X"03",
													6230	=>X"e0",
													6231	=>X"3f",
													6232	=>X"8f",
													6233	=>X"0f",
													6234	=>X"c7",
													6235	=>X"e0",
													6236	=>X"00",
													6237	=>X"00",
													6238	=>X"00",
													6239	=>X"00",
													6240	=>X"00",
													6241	=>X"00",
													6242	=>X"00",
													6243	=>X"00",
													6244	=>X"00",
													6245	=>X"00",
													6246	=>X"00",
													6247	=>X"00",
													6248	=>X"00",
													6249	=>X"00",
													6250	=>X"00",
													6251	=>X"00",
													6252	=>X"00",
													6253	=>X"00",
													6254	=>X"00",
													6255	=>X"00",
													6256	=>X"00",
													6257	=>X"00",
													6258	=>X"00",
													6259	=>X"00",
													6260	=>X"00",
													6261	=>X"00",
													6262	=>X"00",
													6263	=>X"00",
													6264	=>X"00",
													6265	=>X"00",
													6266	=>X"00",
													6267	=>X"00",
													6268	=>X"00",
													6269	=>X"03",
													6270	=>X"f0",
													6271	=>X"1f",
													6272	=>X"ff",
													6273	=>X"7f",
													6274	=>X"87",
													6275	=>X"e0",
													6276	=>X"00",
													6277	=>X"00",
													6278	=>X"00",
													6279	=>X"00",
													6280	=>X"00",
													6281	=>X"00",
													6282	=>X"00",
													6283	=>X"00",
													6284	=>X"00",
													6285	=>X"00",
													6286	=>X"00",
													6287	=>X"00",
													6288	=>X"00",
													6289	=>X"00",
													6290	=>X"00",
													6291	=>X"00",
													6292	=>X"00",
													6293	=>X"00",
													6294	=>X"00",
													6295	=>X"00",
													6296	=>X"00",
													6297	=>X"00",
													6298	=>X"00",
													6299	=>X"00",
													6300	=>X"00",
													6301	=>X"00",
													6302	=>X"00",
													6303	=>X"00",
													6304	=>X"00",
													6305	=>X"00",
													6306	=>X"00",
													6307	=>X"00",
													6308	=>X"00",
													6309	=>X"03",
													6310	=>X"f0",
													6311	=>X"0f",
													6312	=>X"ff",
													6313	=>X"ff",
													6314	=>X"87",
													6315	=>X"c0",
													6316	=>X"00",
													6317	=>X"00",
													6318	=>X"00",
													6319	=>X"00",
													6320	=>X"00",
													6321	=>X"00",
													6322	=>X"00",
													6323	=>X"00",
													6324	=>X"00",
													6325	=>X"00",
													6326	=>X"00",
													6327	=>X"00",
													6328	=>X"00",
													6329	=>X"00",
													6330	=>X"00",
													6331	=>X"00",
													6332	=>X"00",
													6333	=>X"00",
													6334	=>X"00",
													6335	=>X"00",
													6336	=>X"00",
													6337	=>X"00",
													6338	=>X"00",
													6339	=>X"00",
													6340	=>X"00",
													6341	=>X"00",
													6342	=>X"00",
													6343	=>X"00",
													6344	=>X"00",
													6345	=>X"00",
													6346	=>X"00",
													6347	=>X"00",
													6348	=>X"00",
													6349	=>X"03",
													6350	=>X"f0",
													6351	=>X"07",
													6352	=>X"ff",
													6353	=>X"ff",
													6354	=>X"07",
													6355	=>X"c0",
													6356	=>X"00",
													6357	=>X"00",
													6358	=>X"00",
													6359	=>X"00",
													6360	=>X"00",
													6361	=>X"00",
													6362	=>X"00",
													6363	=>X"00",
													6364	=>X"00",
													6365	=>X"00",
													6366	=>X"00",
													6367	=>X"00",
													6368	=>X"00",
													6369	=>X"00",
													6370	=>X"00",
													6371	=>X"00",
													6372	=>X"00",
													6373	=>X"00",
													6374	=>X"00",
													6375	=>X"00",
													6376	=>X"00",
													6377	=>X"00",
													6378	=>X"00",
													6379	=>X"00",
													6380	=>X"00",
													6381	=>X"00",
													6382	=>X"00",
													6383	=>X"00",
													6384	=>X"00",
													6385	=>X"00",
													6386	=>X"00",
													6387	=>X"00",
													6388	=>X"00",
													6389	=>X"03",
													6390	=>X"f0",
													6391	=>X"03",
													6392	=>X"ff",
													6393	=>X"fe",
													6394	=>X"0f",
													6395	=>X"c0",
													6396	=>X"00",
													6397	=>X"00",
													6398	=>X"00",
													6399	=>X"00",
													6400	=>X"00",
													6401	=>X"00",
													6402	=>X"00",
													6403	=>X"00",
													6404	=>X"00",
													6405	=>X"00",
													6406	=>X"00",
													6407	=>X"00",
													6408	=>X"00",
													6409	=>X"00",
													6410	=>X"00",
													6411	=>X"00",
													6412	=>X"00",
													6413	=>X"00",
													6414	=>X"00",
													6415	=>X"00",
													6416	=>X"00",
													6417	=>X"00",
													6418	=>X"00",
													6419	=>X"00",
													6420	=>X"00",
													6421	=>X"00",
													6422	=>X"00",
													6423	=>X"00",
													6424	=>X"00",
													6425	=>X"00",
													6426	=>X"00",
													6427	=>X"00",
													6428	=>X"00",
													6429	=>X"01",
													6430	=>X"f0",
													6431	=>X"01",
													6432	=>X"ff",
													6433	=>X"fc",
													6434	=>X"0f",
													6435	=>X"c0",
													6436	=>X"00",
													6437	=>X"00",
													6438	=>X"00",
													6439	=>X"00",
													6440	=>X"00",
													6441	=>X"00",
													6442	=>X"00",
													6443	=>X"00",
													6444	=>X"00",
													6445	=>X"00",
													6446	=>X"00",
													6447	=>X"00",
													6448	=>X"00",
													6449	=>X"00",
													6450	=>X"00",
													6451	=>X"00",
													6452	=>X"00",
													6453	=>X"00",
													6454	=>X"00",
													6455	=>X"00",
													6456	=>X"00",
													6457	=>X"00",
													6458	=>X"00",
													6459	=>X"00",
													6460	=>X"00",
													6461	=>X"00",
													6462	=>X"00",
													6463	=>X"00",
													6464	=>X"00",
													6465	=>X"00",
													6466	=>X"00",
													6467	=>X"00",
													6468	=>X"00",
													6469	=>X"01",
													6470	=>X"f0",
													6471	=>X"00",
													6472	=>X"3f",
													6473	=>X"e0",
													6474	=>X"0f",
													6475	=>X"c0",
													6476	=>X"00",
													6477	=>X"00",
													6478	=>X"00",
													6479	=>X"00",
													6480	=>X"00",
													6481	=>X"00",
													6482	=>X"00",
													6483	=>X"00",
													6484	=>X"00",
													6485	=>X"00",
													6486	=>X"00",
													6487	=>X"00",
													6488	=>X"00",
													6489	=>X"00",
													6490	=>X"00",
													6491	=>X"00",
													6492	=>X"00",
													6493	=>X"00",
													6494	=>X"00",
													6495	=>X"00",
													6496	=>X"00",
													6497	=>X"00",
													6498	=>X"00",
													6499	=>X"00",
													6500	=>X"00",
													6501	=>X"00",
													6502	=>X"00",
													6503	=>X"00",
													6504	=>X"00",
													6505	=>X"00",
													6506	=>X"00",
													6507	=>X"00",
													6508	=>X"00",
													6509	=>X"01",
													6510	=>X"f8",
													6511	=>X"3c",
													6512	=>X"00",
													6513	=>X"00",
													6514	=>X"0f",
													6515	=>X"80",
													6516	=>X"00",
													6517	=>X"00",
													6518	=>X"00",
													6519	=>X"00",
													6520	=>X"00",
													6521	=>X"00",
													6522	=>X"00",
													6523	=>X"00",
													6524	=>X"00",
													6525	=>X"00",
													6526	=>X"00",
													6527	=>X"00",
													6528	=>X"00",
													6529	=>X"00",
													6530	=>X"00",
													6531	=>X"00",
													6532	=>X"00",
													6533	=>X"00",
													6534	=>X"00",
													6535	=>X"00",
													6536	=>X"00",
													6537	=>X"00",
													6538	=>X"00",
													6539	=>X"00",
													6540	=>X"00",
													6541	=>X"00",
													6542	=>X"00",
													6543	=>X"00",
													6544	=>X"00",
													6545	=>X"00",
													6546	=>X"00",
													6547	=>X"00",
													6548	=>X"00",
													6549	=>X"01",
													6550	=>X"f8",
													6551	=>X"3f",
													6552	=>X"80",
													6553	=>X"00",
													6554	=>X"0f",
													6555	=>X"80",
													6556	=>X"00",
													6557	=>X"00",
													6558	=>X"00",
													6559	=>X"00",
													6560	=>X"00",
													6561	=>X"00",
													6562	=>X"00",
													6563	=>X"00",
													6564	=>X"00",
													6565	=>X"00",
													6566	=>X"00",
													6567	=>X"00",
													6568	=>X"00",
													6569	=>X"00",
													6570	=>X"00",
													6571	=>X"00",
													6572	=>X"00",
													6573	=>X"00",
													6574	=>X"00",
													6575	=>X"00",
													6576	=>X"00",
													6577	=>X"00",
													6578	=>X"00",
													6579	=>X"00",
													6580	=>X"00",
													6581	=>X"00",
													6582	=>X"00",
													6583	=>X"00",
													6584	=>X"00",
													6585	=>X"00",
													6586	=>X"00",
													6587	=>X"00",
													6588	=>X"00",
													6589	=>X"01",
													6590	=>X"f8",
													6591	=>X"3f",
													6592	=>X"e0",
													6593	=>X"00",
													6594	=>X"1f",
													6595	=>X"80",
													6596	=>X"00",
													6597	=>X"00",
													6598	=>X"00",
													6599	=>X"00",
													6600	=>X"00",
													6601	=>X"00",
													6602	=>X"00",
													6603	=>X"00",
													6604	=>X"00",
													6605	=>X"00",
													6606	=>X"00",
													6607	=>X"00",
													6608	=>X"00",
													6609	=>X"00",
													6610	=>X"00",
													6611	=>X"00",
													6612	=>X"00",
													6613	=>X"00",
													6614	=>X"00",
													6615	=>X"00",
													6616	=>X"00",
													6617	=>X"00",
													6618	=>X"00",
													6619	=>X"00",
													6620	=>X"00",
													6621	=>X"00",
													6622	=>X"00",
													6623	=>X"00",
													6624	=>X"00",
													6625	=>X"00",
													6626	=>X"00",
													6627	=>X"00",
													6628	=>X"00",
													6629	=>X"00",
													6630	=>X"f8",
													6631	=>X"3f",
													6632	=>X"f8",
													6633	=>X"00",
													6634	=>X"1f",
													6635	=>X"80",
													6636	=>X"00",
													6637	=>X"00",
													6638	=>X"00",
													6639	=>X"00",
													6640	=>X"00",
													6641	=>X"00",
													6642	=>X"00",
													6643	=>X"00",
													6644	=>X"00",
													6645	=>X"00",
													6646	=>X"00",
													6647	=>X"00",
													6648	=>X"00",
													6649	=>X"00",
													6650	=>X"00",
													6651	=>X"00",
													6652	=>X"00",
													6653	=>X"00",
													6654	=>X"00",
													6655	=>X"00",
													6656	=>X"00",
													6657	=>X"00",
													6658	=>X"00",
													6659	=>X"00",
													6660	=>X"00",
													6661	=>X"00",
													6662	=>X"00",
													6663	=>X"00",
													6664	=>X"00",
													6665	=>X"00",
													6666	=>X"00",
													6667	=>X"00",
													6668	=>X"00",
													6669	=>X"00",
													6670	=>X"fc",
													6671	=>X"1f",
													6672	=>X"fe",
													6673	=>X"00",
													6674	=>X"1f",
													6675	=>X"80",
													6676	=>X"00",
													6677	=>X"00",
													6678	=>X"00",
													6679	=>X"00",
													6680	=>X"00",
													6681	=>X"00",
													6682	=>X"00",
													6683	=>X"00",
													6684	=>X"00",
													6685	=>X"00",
													6686	=>X"00",
													6687	=>X"00",
													6688	=>X"00",
													6689	=>X"00",
													6690	=>X"00",
													6691	=>X"00",
													6692	=>X"00",
													6693	=>X"00",
													6694	=>X"00",
													6695	=>X"00",
													6696	=>X"00",
													6697	=>X"00",
													6698	=>X"00",
													6699	=>X"00",
													6700	=>X"00",
													6701	=>X"00",
													6702	=>X"00",
													6703	=>X"00",
													6704	=>X"00",
													6705	=>X"00",
													6706	=>X"00",
													6707	=>X"00",
													6708	=>X"00",
													6709	=>X"00",
													6710	=>X"fc",
													6711	=>X"18",
													6712	=>X"ff",
													6713	=>X"80",
													6714	=>X"1f",
													6715	=>X"00",
													6716	=>X"00",
													6717	=>X"00",
													6718	=>X"00",
													6719	=>X"00",
													6720	=>X"00",
													6721	=>X"00",
													6722	=>X"00",
													6723	=>X"00",
													6724	=>X"00",
													6725	=>X"00",
													6726	=>X"00",
													6727	=>X"00",
													6728	=>X"00",
													6729	=>X"00",
													6730	=>X"00",
													6731	=>X"00",
													6732	=>X"00",
													6733	=>X"00",
													6734	=>X"00",
													6735	=>X"00",
													6736	=>X"00",
													6737	=>X"00",
													6738	=>X"00",
													6739	=>X"00",
													6740	=>X"00",
													6741	=>X"00",
													6742	=>X"00",
													6743	=>X"00",
													6744	=>X"00",
													6745	=>X"00",
													6746	=>X"00",
													6747	=>X"00",
													6748	=>X"00",
													6749	=>X"00",
													6750	=>X"fc",
													6751	=>X"18",
													6752	=>X"1f",
													6753	=>X"c0",
													6754	=>X"3f",
													6755	=>X"00",
													6756	=>X"00",
													6757	=>X"00",
													6758	=>X"00",
													6759	=>X"00",
													6760	=>X"00",
													6761	=>X"00",
													6762	=>X"00",
													6763	=>X"00",
													6764	=>X"00",
													6765	=>X"00",
													6766	=>X"00",
													6767	=>X"00",
													6768	=>X"00",
													6769	=>X"00",
													6770	=>X"00",
													6771	=>X"00",
													6772	=>X"00",
													6773	=>X"00",
													6774	=>X"00",
													6775	=>X"00",
													6776	=>X"00",
													6777	=>X"00",
													6778	=>X"00",
													6779	=>X"00",
													6780	=>X"00",
													6781	=>X"00",
													6782	=>X"00",
													6783	=>X"00",
													6784	=>X"00",
													6785	=>X"00",
													6786	=>X"00",
													6787	=>X"00",
													6788	=>X"00",
													6789	=>X"00",
													6790	=>X"7c",
													6791	=>X"00",
													6792	=>X"07",
													6793	=>X"e0",
													6794	=>X"3f",
													6795	=>X"00",
													6796	=>X"00",
													6797	=>X"00",
													6798	=>X"00",
													6799	=>X"00",
													6800	=>X"00",
													6801	=>X"00",
													6802	=>X"00",
													6803	=>X"00",
													6804	=>X"00",
													6805	=>X"00",
													6806	=>X"00",
													6807	=>X"00",
													6808	=>X"00",
													6809	=>X"00",
													6810	=>X"00",
													6811	=>X"00",
													6812	=>X"00",
													6813	=>X"00",
													6814	=>X"00",
													6815	=>X"00",
													6816	=>X"00",
													6817	=>X"00",
													6818	=>X"00",
													6819	=>X"00",
													6820	=>X"00",
													6821	=>X"00",
													6822	=>X"00",
													6823	=>X"00",
													6824	=>X"00",
													6825	=>X"00",
													6826	=>X"00",
													6827	=>X"00",
													6828	=>X"00",
													6829	=>X"00",
													6830	=>X"7e",
													6831	=>X"00",
													6832	=>X"01",
													6833	=>X"f0",
													6834	=>X"3f",
													6835	=>X"00",
													6836	=>X"00",
													6837	=>X"00",
													6838	=>X"00",
													6839	=>X"00",
													6840	=>X"00",
													6841	=>X"00",
													6842	=>X"00",
													6843	=>X"00",
													6844	=>X"00",
													6845	=>X"00",
													6846	=>X"00",
													6847	=>X"00",
													6848	=>X"00",
													6849	=>X"00",
													6850	=>X"00",
													6851	=>X"00",
													6852	=>X"00",
													6853	=>X"00",
													6854	=>X"00",
													6855	=>X"00",
													6856	=>X"00",
													6857	=>X"00",
													6858	=>X"00",
													6859	=>X"00",
													6860	=>X"00",
													6861	=>X"00",
													6862	=>X"00",
													6863	=>X"00",
													6864	=>X"00",
													6865	=>X"00",
													6866	=>X"00",
													6867	=>X"00",
													6868	=>X"00",
													6869	=>X"00",
													6870	=>X"7e",
													6871	=>X"00",
													6872	=>X"00",
													6873	=>X"fe",
													6874	=>X"7e",
													6875	=>X"00",
													6876	=>X"00",
													6877	=>X"00",
													6878	=>X"00",
													6879	=>X"00",
													6880	=>X"00",
													6881	=>X"00",
													6882	=>X"00",
													6883	=>X"00",
													6884	=>X"00",
													6885	=>X"00",
													6886	=>X"00",
													6887	=>X"00",
													6888	=>X"00",
													6889	=>X"00",
													6890	=>X"00",
													6891	=>X"00",
													6892	=>X"00",
													6893	=>X"00",
													6894	=>X"00",
													6895	=>X"00",
													6896	=>X"00",
													6897	=>X"00",
													6898	=>X"00",
													6899	=>X"00",
													6900	=>X"00",
													6901	=>X"00",
													6902	=>X"00",
													6903	=>X"00",
													6904	=>X"00",
													6905	=>X"00",
													6906	=>X"00",
													6907	=>X"00",
													6908	=>X"00",
													6909	=>X"00",
													6910	=>X"7e",
													6911	=>X"00",
													6912	=>X"00",
													6913	=>X"7e",
													6914	=>X"7e",
													6915	=>X"00",
													6916	=>X"00",
													6917	=>X"00",
													6918	=>X"00",
													6919	=>X"00",
													6920	=>X"00",
													6921	=>X"00",
													6922	=>X"00",
													6923	=>X"00",
													6924	=>X"00",
													6925	=>X"00",
													6926	=>X"00",
													6927	=>X"00",
													6928	=>X"00",
													6929	=>X"00",
													6930	=>X"00",
													6931	=>X"00",
													6932	=>X"00",
													6933	=>X"00",
													6934	=>X"00",
													6935	=>X"00",
													6936	=>X"00",
													6937	=>X"00",
													6938	=>X"00",
													6939	=>X"00",
													6940	=>X"00",
													6941	=>X"00",
													6942	=>X"00",
													6943	=>X"00",
													6944	=>X"00",
													6945	=>X"00",
													6946	=>X"00",
													6947	=>X"00",
													6948	=>X"00",
													6949	=>X"00",
													6950	=>X"3f",
													6951	=>X"00",
													6952	=>X"00",
													6953	=>X"3e",
													6954	=>X"7e",
													6955	=>X"00",
													6956	=>X"00",
													6957	=>X"00",
													6958	=>X"00",
													6959	=>X"00",
													6960	=>X"00",
													6961	=>X"00",
													6962	=>X"00",
													6963	=>X"00",
													6964	=>X"00",
													6965	=>X"00",
													6966	=>X"00",
													6967	=>X"00",
													6968	=>X"00",
													6969	=>X"00",
													6970	=>X"00",
													6971	=>X"00",
													6972	=>X"00",
													6973	=>X"00",
													6974	=>X"00",
													6975	=>X"00",
													6976	=>X"00",
													6977	=>X"00",
													6978	=>X"00",
													6979	=>X"00",
													6980	=>X"00",
													6981	=>X"00",
													6982	=>X"00",
													6983	=>X"00",
													6984	=>X"00",
													6985	=>X"00",
													6986	=>X"00",
													6987	=>X"00",
													6988	=>X"00",
													6989	=>X"00",
													6990	=>X"3f",
													6991	=>X"06",
													6992	=>X"00",
													6993	=>X"1e",
													6994	=>X"fc",
													6995	=>X"00",
													6996	=>X"00",
													6997	=>X"00",
													6998	=>X"00",
													6999	=>X"00",
													7000	=>X"00",
													7001	=>X"00",
													7002	=>X"00",
													7003	=>X"00",
													7004	=>X"00",
													7005	=>X"00",
													7006	=>X"00",
													7007	=>X"00",
													7008	=>X"00",
													7009	=>X"00",
													7010	=>X"00",
													7011	=>X"00",
													7012	=>X"00",
													7013	=>X"00",
													7014	=>X"00",
													7015	=>X"00",
													7016	=>X"00",
													7017	=>X"00",
													7018	=>X"00",
													7019	=>X"00",
													7020	=>X"00",
													7021	=>X"00",
													7022	=>X"00",
													7023	=>X"00",
													7024	=>X"00",
													7025	=>X"00",
													7026	=>X"00",
													7027	=>X"00",
													7028	=>X"00",
													7029	=>X"00",
													7030	=>X"3f",
													7031	=>X"07",
													7032	=>X"00",
													7033	=>X"1c",
													7034	=>X"fc",
													7035	=>X"00",
													7036	=>X"00",
													7037	=>X"00",
													7038	=>X"00",
													7039	=>X"00",
													7040	=>X"00",
													7041	=>X"00",
													7042	=>X"00",
													7043	=>X"00",
													7044	=>X"00",
													7045	=>X"00",
													7046	=>X"00",
													7047	=>X"00",
													7048	=>X"00",
													7049	=>X"00",
													7050	=>X"00",
													7051	=>X"00",
													7052	=>X"00",
													7053	=>X"00",
													7054	=>X"00",
													7055	=>X"00",
													7056	=>X"00",
													7057	=>X"00",
													7058	=>X"00",
													7059	=>X"00",
													7060	=>X"00",
													7061	=>X"00",
													7062	=>X"00",
													7063	=>X"00",
													7064	=>X"00",
													7065	=>X"00",
													7066	=>X"00",
													7067	=>X"00",
													7068	=>X"00",
													7069	=>X"00",
													7070	=>X"1f",
													7071	=>X"87",
													7072	=>X"e0",
													7073	=>X"1d",
													7074	=>X"fc",
													7075	=>X"00",
													7076	=>X"00",
													7077	=>X"00",
													7078	=>X"00",
													7079	=>X"00",
													7080	=>X"00",
													7081	=>X"00",
													7082	=>X"00",
													7083	=>X"00",
													7084	=>X"00",
													7085	=>X"00",
													7086	=>X"00",
													7087	=>X"00",
													7088	=>X"00",
													7089	=>X"00",
													7090	=>X"00",
													7091	=>X"00",
													7092	=>X"00",
													7093	=>X"00",
													7094	=>X"00",
													7095	=>X"00",
													7096	=>X"00",
													7097	=>X"00",
													7098	=>X"00",
													7099	=>X"00",
													7100	=>X"00",
													7101	=>X"00",
													7102	=>X"00",
													7103	=>X"00",
													7104	=>X"00",
													7105	=>X"00",
													7106	=>X"00",
													7107	=>X"00",
													7108	=>X"00",
													7109	=>X"00",
													7110	=>X"1f",
													7111	=>X"83",
													7112	=>X"fe",
													7113	=>X"3d",
													7114	=>X"f8",
													7115	=>X"00",
													7116	=>X"00",
													7117	=>X"00",
													7118	=>X"00",
													7119	=>X"00",
													7120	=>X"00",
													7121	=>X"00",
													7122	=>X"00",
													7123	=>X"00",
													7124	=>X"00",
													7125	=>X"00",
													7126	=>X"00",
													7127	=>X"00",
													7128	=>X"00",
													7129	=>X"00",
													7130	=>X"00",
													7131	=>X"00",
													7132	=>X"00",
													7133	=>X"00",
													7134	=>X"00",
													7135	=>X"00",
													7136	=>X"00",
													7137	=>X"00",
													7138	=>X"00",
													7139	=>X"00",
													7140	=>X"00",
													7141	=>X"00",
													7142	=>X"00",
													7143	=>X"00",
													7144	=>X"00",
													7145	=>X"00",
													7146	=>X"00",
													7147	=>X"00",
													7148	=>X"00",
													7149	=>X"00",
													7150	=>X"1f",
													7151	=>X"c3",
													7152	=>X"ff",
													7153	=>X"f9",
													7154	=>X"f8",
													7155	=>X"00",
													7156	=>X"00",
													7157	=>X"00",
													7158	=>X"00",
													7159	=>X"00",
													7160	=>X"00",
													7161	=>X"00",
													7162	=>X"00",
													7163	=>X"00",
													7164	=>X"00",
													7165	=>X"00",
													7166	=>X"00",
													7167	=>X"00",
													7168	=>X"00",
													7169	=>X"00",
													7170	=>X"00",
													7171	=>X"00",
													7172	=>X"00",
													7173	=>X"00",
													7174	=>X"00",
													7175	=>X"00",
													7176	=>X"00",
													7177	=>X"00",
													7178	=>X"00",
													7179	=>X"00",
													7180	=>X"00",
													7181	=>X"00",
													7182	=>X"00",
													7183	=>X"00",
													7184	=>X"00",
													7185	=>X"00",
													7186	=>X"00",
													7187	=>X"00",
													7188	=>X"00",
													7189	=>X"00",
													7190	=>X"0f",
													7191	=>X"c1",
													7192	=>X"ff",
													7193	=>X"f3",
													7194	=>X"f8",
													7195	=>X"00",
													7196	=>X"00",
													7197	=>X"00",
													7198	=>X"00",
													7199	=>X"00",
													7200	=>X"00",
													7201	=>X"00",
													7202	=>X"00",
													7203	=>X"00",
													7204	=>X"00",
													7205	=>X"00",
													7206	=>X"00",
													7207	=>X"00",
													7208	=>X"00",
													7209	=>X"00",
													7210	=>X"00",
													7211	=>X"00",
													7212	=>X"00",
													7213	=>X"00",
													7214	=>X"00",
													7215	=>X"00",
													7216	=>X"00",
													7217	=>X"00",
													7218	=>X"00",
													7219	=>X"00",
													7220	=>X"00",
													7221	=>X"00",
													7222	=>X"00",
													7223	=>X"00",
													7224	=>X"00",
													7225	=>X"00",
													7226	=>X"00",
													7227	=>X"00",
													7228	=>X"00",
													7229	=>X"00",
													7230	=>X"0f",
													7231	=>X"c1",
													7232	=>X"ff",
													7233	=>X"f3",
													7234	=>X"f0",
													7235	=>X"00",
													7236	=>X"00",
													7237	=>X"00",
													7238	=>X"00",
													7239	=>X"00",
													7240	=>X"00",
													7241	=>X"00",
													7242	=>X"00",
													7243	=>X"00",
													7244	=>X"00",
													7245	=>X"00",
													7246	=>X"00",
													7247	=>X"00",
													7248	=>X"00",
													7249	=>X"00",
													7250	=>X"00",
													7251	=>X"00",
													7252	=>X"00",
													7253	=>X"00",
													7254	=>X"00",
													7255	=>X"00",
													7256	=>X"00",
													7257	=>X"00",
													7258	=>X"00",
													7259	=>X"00",
													7260	=>X"00",
													7261	=>X"00",
													7262	=>X"00",
													7263	=>X"00",
													7264	=>X"00",
													7265	=>X"00",
													7266	=>X"00",
													7267	=>X"00",
													7268	=>X"00",
													7269	=>X"00",
													7270	=>X"07",
													7271	=>X"e0",
													7272	=>X"df",
													7273	=>X"e7",
													7274	=>X"f0",
													7275	=>X"00",
													7276	=>X"00",
													7277	=>X"00",
													7278	=>X"00",
													7279	=>X"00",
													7280	=>X"00",
													7281	=>X"00",
													7282	=>X"00",
													7283	=>X"00",
													7284	=>X"00",
													7285	=>X"00",
													7286	=>X"00",
													7287	=>X"00",
													7288	=>X"00",
													7289	=>X"00",
													7290	=>X"00",
													7291	=>X"00",
													7292	=>X"00",
													7293	=>X"00",
													7294	=>X"00",
													7295	=>X"00",
													7296	=>X"00",
													7297	=>X"00",
													7298	=>X"00",
													7299	=>X"00",
													7300	=>X"00",
													7301	=>X"00",
													7302	=>X"00",
													7303	=>X"00",
													7304	=>X"00",
													7305	=>X"00",
													7306	=>X"00",
													7307	=>X"00",
													7308	=>X"00",
													7309	=>X"00",
													7310	=>X"07",
													7311	=>X"f0",
													7312	=>X"c1",
													7313	=>X"ef",
													7314	=>X"e0",
													7315	=>X"00",
													7316	=>X"00",
													7317	=>X"00",
													7318	=>X"00",
													7319	=>X"00",
													7320	=>X"00",
													7321	=>X"00",
													7322	=>X"00",
													7323	=>X"00",
													7324	=>X"00",
													7325	=>X"00",
													7326	=>X"00",
													7327	=>X"00",
													7328	=>X"00",
													7329	=>X"00",
													7330	=>X"00",
													7331	=>X"00",
													7332	=>X"00",
													7333	=>X"00",
													7334	=>X"00",
													7335	=>X"00",
													7336	=>X"00",
													7337	=>X"00",
													7338	=>X"00",
													7339	=>X"00",
													7340	=>X"00",
													7341	=>X"00",
													7342	=>X"00",
													7343	=>X"00",
													7344	=>X"00",
													7345	=>X"00",
													7346	=>X"00",
													7347	=>X"00",
													7348	=>X"00",
													7349	=>X"00",
													7350	=>X"07",
													7351	=>X"f0",
													7352	=>X"00",
													7353	=>X"ef",
													7354	=>X"e0",
													7355	=>X"00",
													7356	=>X"00",
													7357	=>X"00",
													7358	=>X"00",
													7359	=>X"00",
													7360	=>X"00",
													7361	=>X"00",
													7362	=>X"00",
													7363	=>X"00",
													7364	=>X"00",
													7365	=>X"00",
													7366	=>X"00",
													7367	=>X"00",
													7368	=>X"00",
													7369	=>X"00",
													7370	=>X"00",
													7371	=>X"00",
													7372	=>X"00",
													7373	=>X"00",
													7374	=>X"00",
													7375	=>X"00",
													7376	=>X"00",
													7377	=>X"00",
													7378	=>X"00",
													7379	=>X"00",
													7380	=>X"00",
													7381	=>X"00",
													7382	=>X"00",
													7383	=>X"00",
													7384	=>X"00",
													7385	=>X"00",
													7386	=>X"00",
													7387	=>X"00",
													7388	=>X"00",
													7389	=>X"00",
													7390	=>X"03",
													7391	=>X"f8",
													7392	=>X"00",
													7393	=>X"9f",
													7394	=>X"c0",
													7395	=>X"00",
													7396	=>X"00",
													7397	=>X"00",
													7398	=>X"00",
													7399	=>X"00",
													7400	=>X"00",
													7401	=>X"00",
													7402	=>X"00",
													7403	=>X"00",
													7404	=>X"00",
													7405	=>X"00",
													7406	=>X"00",
													7407	=>X"00",
													7408	=>X"00",
													7409	=>X"00",
													7410	=>X"00",
													7411	=>X"00",
													7412	=>X"00",
													7413	=>X"00",
													7414	=>X"00",
													7415	=>X"00",
													7416	=>X"00",
													7417	=>X"00",
													7418	=>X"00",
													7419	=>X"00",
													7420	=>X"00",
													7421	=>X"00",
													7422	=>X"00",
													7423	=>X"00",
													7424	=>X"00",
													7425	=>X"00",
													7426	=>X"00",
													7427	=>X"00",
													7428	=>X"00",
													7429	=>X"00",
													7430	=>X"03",
													7431	=>X"f8",
													7432	=>X"00",
													7433	=>X"1f",
													7434	=>X"c0",
													7435	=>X"00",
													7436	=>X"00",
													7437	=>X"00",
													7438	=>X"00",
													7439	=>X"00",
													7440	=>X"00",
													7441	=>X"00",
													7442	=>X"00",
													7443	=>X"00",
													7444	=>X"00",
													7445	=>X"00",
													7446	=>X"00",
													7447	=>X"00",
													7448	=>X"00",
													7449	=>X"00",
													7450	=>X"00",
													7451	=>X"00",
													7452	=>X"00",
													7453	=>X"00",
													7454	=>X"00",
													7455	=>X"00",
													7456	=>X"00",
													7457	=>X"00",
													7458	=>X"00",
													7459	=>X"00",
													7460	=>X"00",
													7461	=>X"00",
													7462	=>X"00",
													7463	=>X"00",
													7464	=>X"00",
													7465	=>X"00",
													7466	=>X"00",
													7467	=>X"00",
													7468	=>X"00",
													7469	=>X"00",
													7470	=>X"01",
													7471	=>X"ff",
													7472	=>X"ff",
													7473	=>X"ff",
													7474	=>X"c0",
													7475	=>X"00",
													7476	=>X"00",
													7477	=>X"00",
													7478	=>X"00",
													7479	=>X"00",
													7480	=>X"00",
													7481	=>X"00",
													7482	=>X"00",
													7483	=>X"00",
													7484	=>X"00",
													7485	=>X"00",
													7486	=>X"00",
													7487	=>X"00",
													7488	=>X"00",
													7489	=>X"00",
													7490	=>X"00",
													7491	=>X"00",
													7492	=>X"00",
													7493	=>X"00",
													7494	=>X"00",
													7495	=>X"00",
													7496	=>X"00",
													7497	=>X"00",
													7498	=>X"00",
													7499	=>X"00",
													7500	=>X"00",
													7501	=>X"00",
													7502	=>X"00",
													7503	=>X"00",
													7504	=>X"00",
													7505	=>X"00",
													7506	=>X"00",
													7507	=>X"00",
													7508	=>X"00",
													7509	=>X"00",
													7510	=>X"01",
													7511	=>X"ff",
													7512	=>X"ff",
													7513	=>X"ff",
													7514	=>X"80",
													7515	=>X"00",
													7516	=>X"00",
													7517	=>X"00",
													7518	=>X"00",
													7519	=>X"00",
													7520	=>X"00",
													7521	=>X"00",
													7522	=>X"00",
													7523	=>X"00",
													7524	=>X"00",
													7525	=>X"00",
													7526	=>X"00",
													7527	=>X"00",
													7528	=>X"00",
													7529	=>X"00",
													7530	=>X"00",
													7531	=>X"00",
													7532	=>X"00",
													7533	=>X"00",
													7534	=>X"00",
													7535	=>X"00",
													7536	=>X"00",
													7537	=>X"00",
													7538	=>X"00",
													7539	=>X"00",
													7540	=>X"00",
													7541	=>X"00",
													7542	=>X"00",
													7543	=>X"00",
													7544	=>X"00",
													7545	=>X"00",
													7546	=>X"00",
													7547	=>X"00",
													7548	=>X"00",
													7549	=>X"00",
													7550	=>X"00",
													7551	=>X"ff",
													7552	=>X"ff",
													7553	=>X"ff",
													7554	=>X"80",
													7555	=>X"00",
													7556	=>X"00",
													7557	=>X"00",
													7558	=>X"00",
													7559	=>X"00",
													7560	=>X"00",
													7561	=>X"00",
													7562	=>X"00",
													7563	=>X"00",
													7564	=>X"00",
													7565	=>X"00",
													7566	=>X"00",
													7567	=>X"00",
													7568	=>X"00",
													7569	=>X"00",
													7570	=>X"00",
													7571	=>X"00",
													7572	=>X"00",
													7573	=>X"00",
													7574	=>X"00",
													7575	=>X"00",
													7576	=>X"00",
													7577	=>X"00",
													7578	=>X"00",
													7579	=>X"00",
													7580	=>X"00",
													7581	=>X"00",
													7582	=>X"00",
													7583	=>X"00",
													7584	=>X"00",
													7585	=>X"00",
													7586	=>X"00",
													7587	=>X"00",
													7588	=>X"00",
													7589	=>X"00",
													7590	=>X"00",
													7591	=>X"ff",
													7592	=>X"ff",
													7593	=>X"ff",
													7594	=>X"00",
													7595	=>X"00",
													7596	=>X"00",
													7597	=>X"00",
													7598	=>X"00",
													7599	=>X"00",
													7600	=>X"00",
													7601	=>X"00",
													7602	=>X"00",
													7603	=>X"00",
													7604	=>X"00",
													7605	=>X"00",
													7606	=>X"00",
													7607	=>X"00",
													7608	=>X"00",
													7609	=>X"00",
													7610	=>X"00",
													7611	=>X"00",
													7612	=>X"00",
													7613	=>X"00",
													7614	=>X"00",
													7615	=>X"00",
													7616	=>X"00",
													7617	=>X"00",
													7618	=>X"00",
													7619	=>X"00",
													7620	=>X"00",
													7621	=>X"00",
													7622	=>X"00",
													7623	=>X"00",
													7624	=>X"00",
													7625	=>X"00",
													7626	=>X"00",
													7627	=>X"00",
													7628	=>X"00",
													7629	=>X"00",
													7630	=>X"00",
													7631	=>X"7f",
													7632	=>X"ff",
													7633	=>X"fe",
													7634	=>X"00",
													7635	=>X"00",
													7636	=>X"00",
													7637	=>X"00",
													7638	=>X"00",
													7639	=>X"00",
													7640	=>X"00",
													7641	=>X"00",
													7642	=>X"00",
													7643	=>X"00",
													7644	=>X"00",
													7645	=>X"00",
													7646	=>X"00",
													7647	=>X"00",
													7648	=>X"00",
													7649	=>X"00",
													7650	=>X"00",
													7651	=>X"00",
													7652	=>X"00",
													7653	=>X"00",
													7654	=>X"00",
													7655	=>X"00",
													7656	=>X"00",
													7657	=>X"00",
													7658	=>X"00",
													7659	=>X"00",
													7660	=>X"00",
													7661	=>X"00",
													7662	=>X"00",
													7663	=>X"00",
													7664	=>X"00",
													7665	=>X"00",
													7666	=>X"00",
													7667	=>X"00",
													7668	=>X"00",
													7669	=>X"00",
													7670	=>X"00",
													7671	=>X"7f",
													7672	=>X"ff",
													7673	=>X"fe",
													7674	=>X"00",
													7675	=>X"00",
													7676	=>X"00",
													7677	=>X"00",
													7678	=>X"00",
													7679	=>X"00",
													7680	=>X"00",
													7681	=>X"00",
													7682	=>X"00",
													7683	=>X"00",
													7684	=>X"00",
													7685	=>X"00",
													7686	=>X"00",
													7687	=>X"00",
													7688	=>X"00",
													7689	=>X"00",
													7690	=>X"00",
													7691	=>X"00",
													7692	=>X"00",
													7693	=>X"00",
													7694	=>X"00",
													7695	=>X"00",
													7696	=>X"00",
													7697	=>X"00",
													7698	=>X"00",
													7699	=>X"00",
													7700	=>X"00",
													7701	=>X"00",
													7702	=>X"00",
													7703	=>X"00",
													7704	=>X"00",
													7705	=>X"00",
													7706	=>X"00",
													7707	=>X"00",
													7708	=>X"00",
													7709	=>X"00",
													7710	=>X"00",
													7711	=>X"3f",
													7712	=>X"ff",
													7713	=>X"fc",
													7714	=>X"00",
													7715	=>X"00",
													7716	=>X"00",
													7717	=>X"00",
													7718	=>X"00",
													7719	=>X"00",
													7720	=>X"00",
													7721	=>X"00",
													7722	=>X"00",
													7723	=>X"00",
													7724	=>X"00",
													7725	=>X"00",
													7726	=>X"00",
													7727	=>X"00",
													7728	=>X"00",
													7729	=>X"00",
													7730	=>X"00",
													7731	=>X"00",
													7732	=>X"00",
													7733	=>X"00",
													7734	=>X"00",
													7735	=>X"00",
													7736	=>X"00",
													7737	=>X"00",
													7738	=>X"00",
													7739	=>X"00",
													7740	=>X"00",
													7741	=>X"00",
													7742	=>X"00",
													7743	=>X"00",
													7744	=>X"00",
													7745	=>X"00",
													7746	=>X"00",
													7747	=>X"00",
													7748	=>X"00",
													7749	=>X"00",
													7750	=>X"00",
													7751	=>X"1f",
													7752	=>X"ff",
													7753	=>X"f8",
													7754	=>X"00",
													7755	=>X"00",
													7756	=>X"00",
													7757	=>X"00",
													7758	=>X"00",
													7759	=>X"00",
													7760	=>X"00",
													7761	=>X"00",
													7762	=>X"00",
													7763	=>X"00",
													7764	=>X"00",
													7765	=>X"00",
													7766	=>X"00",
													7767	=>X"00",
													7768	=>X"00",
													7769	=>X"00",
													7770	=>X"00",
													7771	=>X"00",
													7772	=>X"00",
													7773	=>X"00",
													7774	=>X"00",
													7775	=>X"00",
													7776	=>X"00",
													7777	=>X"00",
													7778	=>X"00",
													7779	=>X"00",
													7780	=>X"00",
													7781	=>X"00",
													7782	=>X"00",
													7783	=>X"00",
													7784	=>X"00",
													7785	=>X"00",
													7786	=>X"00",
													7787	=>X"00",
													7788	=>X"00",
													7789	=>X"00",
													7790	=>X"00",
													7791	=>X"0f",
													7792	=>X"ff",
													7793	=>X"f0",
													7794	=>X"00",
													7795	=>X"00",
													7796	=>X"00",
													7797	=>X"00",
													7798	=>X"00",
													7799	=>X"00",
													7800	=>X"00",
													7801	=>X"00",
													7802	=>X"00",
													7803	=>X"00",
													7804	=>X"00",
													7805	=>X"00",
													7806	=>X"00",
													7807	=>X"00",
													7808	=>X"00",
													7809	=>X"00",
													7810	=>X"00",
													7811	=>X"00",
													7812	=>X"00",
													7813	=>X"00",
													7814	=>X"00",
													7815	=>X"00",
													7816	=>X"00",
													7817	=>X"00",
													7818	=>X"00",
													7819	=>X"00",
													7820	=>X"00",
													7821	=>X"00",
													7822	=>X"00",
													7823	=>X"00",
													7824	=>X"00",
													7825	=>X"00",
													7826	=>X"00",
													7827	=>X"00",
													7828	=>X"00",
													7829	=>X"00",
													7830	=>X"00",
													7831	=>X"00",
													7832	=>X"00",
													7833	=>X"00",
													7834	=>X"00",
													7835	=>X"00",
													7836	=>X"00",
													7837	=>X"00",
													7838	=>X"00",
													7839	=>X"00",
													7840	=>X"00",
													7841	=>X"00",
													7842	=>X"00",
													7843	=>X"00",
													7844	=>X"00",
													7845	=>X"00",
													7846	=>X"00",
													7847	=>X"00",
													7848	=>X"00",
													7849	=>X"00",
													7850	=>X"00",
													7851	=>X"00",
													7852	=>X"00",
													7853	=>X"00",
													7854	=>X"00",
													7855	=>X"00",
													7856	=>X"00",
													7857	=>X"00",
													7858	=>X"00",
													7859	=>X"00",
													7860	=>X"00",
													7861	=>X"00",
													7862	=>X"00",
													7863	=>X"00",
													7864	=>X"00",
													7865	=>X"00",
													7866	=>X"00",
													7867	=>X"00",
													7868	=>X"00",
													7869	=>X"00",
													7870	=>X"00",
													7871	=>X"00",
													7872	=>X"00",
													7873	=>X"00",
													7874	=>X"00",
													7875	=>X"00",
													7876	=>X"00",
													7877	=>X"00",
													7878	=>X"00",
													7879	=>X"00",
													7880	=>X"00",
													7881	=>X"00",
													7882	=>X"00",
													7883	=>X"00",
													7884	=>X"00",
													7885	=>X"00",
													7886	=>X"00",
													7887	=>X"00",
													7888	=>X"00",
													7889	=>X"00",
													7890	=>X"00",
													7891	=>X"00",
													7892	=>X"00",
													7893	=>X"00",
													7894	=>X"00",
													7895	=>X"00",
													7896	=>X"00",
													7897	=>X"00",
													7898	=>X"00",
													7899	=>X"00",
													7900	=>X"00",
													7901	=>X"00",
													7902	=>X"00",
													7903	=>X"00",
													7904	=>X"00",
													7905	=>X"00",
													7906	=>X"00",
													7907	=>X"00",
													7908	=>X"00",
													7909	=>X"00",
													7910	=>X"00",
													7911	=>X"00",
													7912	=>X"00",
													7913	=>X"00",
													7914	=>X"00",
													7915	=>X"00",
													7916	=>X"00",
													7917	=>X"00",
													7918	=>X"00",
													7919	=>X"00",
													7920	=>X"00",
													7921	=>X"00",
													7922	=>X"00",
													7923	=>X"00",
													7924	=>X"00",
													7925	=>X"00",
													7926	=>X"00",
													7927	=>X"00",
													7928	=>X"00",
													7929	=>X"00",
													7930	=>X"00",
													7931	=>X"00",
													7932	=>X"00",
													7933	=>X"00",
													7934	=>X"00",
													7935	=>X"00",
													7936	=>X"00",
													7937	=>X"00",
													7938	=>X"00",
													7939	=>X"00",
													7940	=>X"00",
													7941	=>X"00",
													7942	=>X"00",
													7943	=>X"00",
													7944	=>X"00",
													7945	=>X"00",
													7946	=>X"00",
													7947	=>X"00",
													7948	=>X"00",
													7949	=>X"00",
													7950	=>X"00",
													7951	=>X"00",
													7952	=>X"00",
													7953	=>X"00",
													7954	=>X"00",
													7955	=>X"00",
													7956	=>X"00",
													7957	=>X"00",
													7958	=>X"00",
													7959	=>X"00",
													7960	=>X"00",
													7961	=>X"00",
													7962	=>X"00",
													7963	=>X"00",
													7964	=>X"00",
													7965	=>X"00",
													7966	=>X"00",
													7967	=>X"00",
													7968	=>X"00",
													7969	=>X"00",
													7970	=>X"00",
													7971	=>X"00",
													7972	=>X"00",
													7973	=>X"00",
													7974	=>X"00",
													7975	=>X"00",
													7976	=>X"00",
													7977	=>X"00",
													7978	=>X"00",
													7979	=>X"00",
													7980	=>X"00",
													7981	=>X"00",
													7982	=>X"00",
													7983	=>X"00",
													7984	=>X"00",
													7985	=>X"00",
													7986	=>X"00",
													7987	=>X"00",
													7988	=>X"00",
													7989	=>X"00",
													7990	=>X"00",
													7991	=>X"00",
													7992	=>X"00",
													7993	=>X"00",
													7994	=>X"00",
													7995	=>X"00",
													7996	=>X"00",
													7997	=>X"00",
													7998	=>X"00",
													7999	=>X"00",
													8000	=>X"00",
													8001	=>X"00",
													8002	=>X"00",
													8003	=>X"00",
													8004	=>X"00",
													8005	=>X"00",
													8006	=>X"00",
													8007	=>X"00",
													8008	=>X"00",
													8009	=>X"00",
													8010	=>X"00",
													8011	=>X"00",
													8012	=>X"00",
													8013	=>X"00",
													8014	=>X"00",
													8015	=>X"00",
													8016	=>X"00",
													8017	=>X"00",
													8018	=>X"00",
													8019	=>X"00",
													8020	=>X"00",
													8021	=>X"00",
													8022	=>X"00",
													8023	=>X"00",
													8024	=>X"00",
													8025	=>X"00",
													8026	=>X"00",
													8027	=>X"00",
													8028	=>X"00",
													8029	=>X"00",
													8030	=>X"00",
													8031	=>X"00",
													8032	=>X"00",
													8033	=>X"00",
													8034	=>X"00",
													8035	=>X"00",
													8036	=>X"00",
													8037	=>X"00",
													8038	=>X"00",
													8039	=>X"00",
													8040	=>X"00",
													8041	=>X"00",
													8042	=>X"00",
													8043	=>X"00",
													8044	=>X"00",
													8045	=>X"00",
													8046	=>X"00",
													8047	=>X"00",
													8048	=>X"00",
													8049	=>X"00",
													8050	=>X"00",
													8051	=>X"00",
													8052	=>X"00",
													8053	=>X"00",
													8054	=>X"00",
													8055	=>X"00",
													8056	=>X"00",
													8057	=>X"00",
													8058	=>X"00",
													8059	=>X"00",
													8060	=>X"00",
													8061	=>X"00",
													8062	=>X"00",
													8063	=>X"00",
													8064	=>X"00",
													8065	=>X"00",
													8066	=>X"00",
													8067	=>X"00",
													8068	=>X"00",
													8069	=>X"00",
													8070	=>X"00",
													8071	=>X"00",
													8072	=>X"00",
													8073	=>X"00",
													8074	=>X"00",
													8075	=>X"00",
													8076	=>X"00",
													8077	=>X"00",
													8078	=>X"00",
													8079	=>X"00",
													8080	=>X"00",
													8081	=>X"00",
													8082	=>X"00",
													8083	=>X"00",
													8084	=>X"00",
													8085	=>X"00",
													8086	=>X"00",
													8087	=>X"00",
													8088	=>X"00",
													8089	=>X"00",
													8090	=>X"00",
													8091	=>X"00",
													8092	=>X"00",
													8093	=>X"00",
													8094	=>X"00",
													8095	=>X"00",
													8096	=>X"00",
													8097	=>X"00",
													8098	=>X"00",
													8099	=>X"00",
													8100	=>X"00",
													8101	=>X"00",
													8102	=>X"00",
													8103	=>X"00",
													8104	=>X"00",
													8105	=>X"00",
													8106	=>X"00",
													8107	=>X"00",
													8108	=>X"00",
													8109	=>X"00",
													8110	=>X"00",
													8111	=>X"00",
													8112	=>X"00",
													8113	=>X"00",
													8114	=>X"00",
													8115	=>X"00",
													8116	=>X"00",
													8117	=>X"00",
													8118	=>X"00",
													8119	=>X"00",
													8120	=>X"00",
													8121	=>X"00",
													8122	=>X"00",
													8123	=>X"00",
													8124	=>X"00",
													8125	=>X"00",
													8126	=>X"00",
													8127	=>X"00",
													8128	=>X"00",
													8129	=>X"00",
													8130	=>X"00",
													8131	=>X"00",
													8132	=>X"00",
													8133	=>X"00",
													8134	=>X"00",
													8135	=>X"00",
													8136	=>X"00",
													8137	=>X"00",
													8138	=>X"00",
													8139	=>X"00",
													8140	=>X"00",
													8141	=>X"00",
													8142	=>X"00",
													8143	=>X"00",
													8144	=>X"00",
													8145	=>X"00",
													8146	=>X"00",
													8147	=>X"00",
													8148	=>X"00",
													8149	=>X"00",
													8150	=>X"00",
													8151	=>X"00",
													8152	=>X"00",
													8153	=>X"00",
													8154	=>X"00",
													8155	=>X"00",
													8156	=>X"00",
													8157	=>X"00",
													8158	=>X"00",
													8159	=>X"00",
													8160	=>X"00",
													8161	=>X"00",
													8162	=>X"00",
													8163	=>X"00",
													8164	=>X"00",
													8165	=>X"00",
													8166	=>X"00",
													8167	=>X"00",
													8168	=>X"00",
													8169	=>X"00",
													8170	=>X"00",
													8171	=>X"00",
													8172	=>X"00",
													8173	=>X"00",
													8174	=>X"00",
													8175	=>X"00",
													8176	=>X"00",
													8177	=>X"00",
													8178	=>X"00",
													8179	=>X"00",
													8180	=>X"00",
													8181	=>X"00",
													8182	=>X"00",
													8183	=>X"00",
													8184	=>X"00",
													8185	=>X"00",
													8186	=>X"00",
													8187	=>X"00",
													8188	=>X"00",
													8189	=>X"00",
													8190	=>X"00",
													8191	=>X"00",
													8192	=>X"00",
													8193	=>X"00",
													8194	=>X"00",
													8195	=>X"00",
													8196	=>X"00",
													8197	=>X"00",
													8198	=>X"00",
													8199	=>X"00",
													8200	=>X"00",
													8201	=>X"00",
													8202	=>X"00",
													8203	=>X"00",
													8204	=>X"00",
													8205	=>X"00",
													8206	=>X"00",
													8207	=>X"00",
													8208	=>X"00",
													8209	=>X"00",
													8210	=>X"00",
													8211	=>X"00",
													8212	=>X"00",
													8213	=>X"00",
													8214	=>X"00",
													8215	=>X"00",
													8216	=>X"00",
													8217	=>X"00",
													8218	=>X"00",
													8219	=>X"00",
													8220	=>X"00",
													8221	=>X"00",
													8222	=>X"00",
													8223	=>X"00",
													8224	=>X"00",
													8225	=>X"00",
													8226	=>X"00",
													8227	=>X"00",
													8228	=>X"00",
													8229	=>X"00",
													8230	=>X"00",
													8231	=>X"00",
													8232	=>X"00",
													8233	=>X"00",
													8234	=>X"00",
													8235	=>X"00",
													8236	=>X"00",
													8237	=>X"00",
													8238	=>X"00",
													8239	=>X"00",
													8240	=>X"00",
													8241	=>X"00",
													8242	=>X"00",
													8243	=>X"00",
													8244	=>X"00",
													8245	=>X"00",
													8246	=>X"00",
													8247	=>X"00",
													8248	=>X"00",
													8249	=>X"00",
													8250	=>X"00",
													8251	=>X"00",
													8252	=>X"00",
													8253	=>X"00",
													8254	=>X"00",
													8255	=>X"00",
													8256	=>X"00",
													8257	=>X"00",
													8258	=>X"00",
													8259	=>X"00",
													8260	=>X"00",
													8261	=>X"00",
													8262	=>X"00",
													8263	=>X"00",
													8264	=>X"00",
													8265	=>X"00",
													8266	=>X"00",
													8267	=>X"00",
													8268	=>X"00",
													8269	=>X"00",
													8270	=>X"00",
													8271	=>X"00",
													8272	=>X"00",
													8273	=>X"00",
													8274	=>X"00",
													8275	=>X"00",
													8276	=>X"00",
													8277	=>X"00",
													8278	=>X"00",
													8279	=>X"00",
													8280	=>X"00",
													8281	=>X"00",
													8282	=>X"00",
													8283	=>X"00",
													8284	=>X"00",
													8285	=>X"00",
													8286	=>X"00",
													8287	=>X"00",
													8288	=>X"00",
													8289	=>X"00",
													8290	=>X"00",
													8291	=>X"00",
													8292	=>X"00",
													8293	=>X"00",
													8294	=>X"00",
													8295	=>X"00",
													8296	=>X"00",
													8297	=>X"00",
													8298	=>X"00",
													8299	=>X"00",
													8300	=>X"00",
													8301	=>X"00",
													8302	=>X"00",
													8303	=>X"00",
													8304	=>X"00",
													8305	=>X"00",
													8306	=>X"00",
													8307	=>X"00",
													8308	=>X"00",
													8309	=>X"00",
													8310	=>X"00",
													8311	=>X"00",
													8312	=>X"00",
													8313	=>X"00",
													8314	=>X"00",
													8315	=>X"00",
													8316	=>X"00",
													8317	=>X"00",
													8318	=>X"00",
													8319	=>X"00",
													8320	=>X"00",
													8321	=>X"00",
													8322	=>X"00",
													8323	=>X"00",
													8324	=>X"00",
													8325	=>X"00",
													8326	=>X"00",
													8327	=>X"00",
													8328	=>X"00",
													8329	=>X"00",
													8330	=>X"00",
													8331	=>X"00",
													8332	=>X"00",
													8333	=>X"00",
													8334	=>X"00",
													8335	=>X"00",
													8336	=>X"00",
													8337	=>X"00",
													8338	=>X"00",
													8339	=>X"00",
													8340	=>X"00",
													8341	=>X"00",
													8342	=>X"00",
													8343	=>X"00",
													8344	=>X"00",
													8345	=>X"00",
													8346	=>X"00",
													8347	=>X"00",
													8348	=>X"00",
													8349	=>X"00",
													8350	=>X"00",
													8351	=>X"00",
													8352	=>X"00",
													8353	=>X"00",
													8354	=>X"00",
													8355	=>X"00",
													8356	=>X"00",
													8357	=>X"00",
													8358	=>X"00",
													8359	=>X"00",
													8360	=>X"00",
													8361	=>X"00",
													8362	=>X"00",
													8363	=>X"00",
													8364	=>X"00",
													8365	=>X"00",
													8366	=>X"00",
													8367	=>X"00",
													8368	=>X"00",
													8369	=>X"00",
													8370	=>X"00",
													8371	=>X"00",
													8372	=>X"00",
													8373	=>X"00",
													8374	=>X"00",
													8375	=>X"00",
													8376	=>X"00",
													8377	=>X"00",
													8378	=>X"00",
													8379	=>X"00",
													8380	=>X"00",
													8381	=>X"00",
													8382	=>X"00",
													8383	=>X"00",
													8384	=>X"00",
													8385	=>X"00",
													8386	=>X"00",
													8387	=>X"00",
													8388	=>X"00",
													8389	=>X"00",
													8390	=>X"00",
													8391	=>X"00",
													8392	=>X"00",
													8393	=>X"00",
													8394	=>X"00",
													8395	=>X"00",
													8396	=>X"00",
													8397	=>X"00",
													8398	=>X"00",
													8399	=>X"00",
													8400	=>X"00",
													8401	=>X"00",
													8402	=>X"00",
													8403	=>X"00",
													8404	=>X"00",
													8405	=>X"00",
													8406	=>X"00",
													8407	=>X"00",
													8408	=>X"00",
													8409	=>X"00",
													8410	=>X"00",
													8411	=>X"00",
													8412	=>X"00",
													8413	=>X"00",
													8414	=>X"00",
													8415	=>X"00",
													8416	=>X"00",
													8417	=>X"00",
													8418	=>X"00",
													8419	=>X"00",
													8420	=>X"00",
													8421	=>X"00",
													8422	=>X"00",
													8423	=>X"00",
													8424	=>X"00",
													8425	=>X"00",
													8426	=>X"00",
													8427	=>X"00",
													8428	=>X"00",
													8429	=>X"00",
													8430	=>X"00",
													8431	=>X"00",
													8432	=>X"00",
													8433	=>X"00",
													8434	=>X"00",
													8435	=>X"00",
													8436	=>X"00",
													8437	=>X"00",
													8438	=>X"00",
													8439	=>X"00",
													8440	=>X"00",
													8441	=>X"00",
													8442	=>X"00",
													8443	=>X"00",
													8444	=>X"00",
													8445	=>X"00",
													8446	=>X"00",
													8447	=>X"00",
													8448	=>X"00",
													8449	=>X"00",
													8450	=>X"00",
													8451	=>X"00",
													8452	=>X"00",
													8453	=>X"00",
													8454	=>X"00",
													8455	=>X"00",
													8456	=>X"00",
													8457	=>X"00",
													8458	=>X"00",
													8459	=>X"00",
													8460	=>X"00",
													8461	=>X"00",
													8462	=>X"00",
													8463	=>X"00",
													8464	=>X"00",
													8465	=>X"00",
													8466	=>X"00",
													8467	=>X"00",
													8468	=>X"00",
													8469	=>X"00",
													8470	=>X"00",
													8471	=>X"00",
													8472	=>X"00",
													8473	=>X"00",
													8474	=>X"00",
													8475	=>X"00",
													8476	=>X"00",
													8477	=>X"00",
													8478	=>X"00",
													8479	=>X"00",
													8480	=>X"00",
													8481	=>X"00",
													8482	=>X"00",
													8483	=>X"00",
													8484	=>X"00",
													8485	=>X"00",
													8486	=>X"00",
													8487	=>X"00",
													8488	=>X"00",
													8489	=>X"00",
													8490	=>X"00",
													8491	=>X"00",
													8492	=>X"00",
													8493	=>X"00",
													8494	=>X"00",
													8495	=>X"00",
													8496	=>X"00",
													8497	=>X"00",
													8498	=>X"00",
													8499	=>X"00",
													8500	=>X"00",
													8501	=>X"00",
													8502	=>X"00",
													8503	=>X"00",
													8504	=>X"00",
													8505	=>X"00",
													8506	=>X"00",
													8507	=>X"00",
													8508	=>X"00",
													8509	=>X"00",
													8510	=>X"00",
													8511	=>X"00",
													8512	=>X"00",
													8513	=>X"00",
													8514	=>X"00",
													8515	=>X"00",
													8516	=>X"00",
													8517	=>X"00",
													8518	=>X"00",
													8519	=>X"00",
													8520	=>X"00",
													8521	=>X"00",
													8522	=>X"00",
													8523	=>X"00",
													8524	=>X"00",
													8525	=>X"00",
													8526	=>X"00",
													8527	=>X"00",
													8528	=>X"00",
													8529	=>X"00",
													8530	=>X"00",
													8531	=>X"00",
													8532	=>X"00",
													8533	=>X"00",
													8534	=>X"00",
													8535	=>X"00",
													8536	=>X"00",
													8537	=>X"00",
													8538	=>X"00",
													8539	=>X"00",
													8540	=>X"00",
													8541	=>X"00",
													8542	=>X"00",
													8543	=>X"00",
													8544	=>X"00",
													8545	=>X"00",
													8546	=>X"00",
													8547	=>X"00",
													8548	=>X"00",
													8549	=>X"00",
													8550	=>X"00",
													8551	=>X"00",
													8552	=>X"00",
													8553	=>X"00",
													8554	=>X"00",
													8555	=>X"00",
													8556	=>X"00",
													8557	=>X"00",
													8558	=>X"00",
													8559	=>X"00",
													8560	=>X"00",
													8561	=>X"00",
													8562	=>X"00",
													8563	=>X"00",
													8564	=>X"00",
													8565	=>X"00",
													8566	=>X"00",
													8567	=>X"00",
													8568	=>X"00",
													8569	=>X"00",
													8570	=>X"00",
													8571	=>X"00",
													8572	=>X"00",
													8573	=>X"00",
													8574	=>X"00",
													8575	=>X"00",
													8576	=>X"00",
													8577	=>X"00",
													8578	=>X"00",
													8579	=>X"00",
													8580	=>X"00",
													8581	=>X"00",
													8582	=>X"00",
													8583	=>X"00",
													8584	=>X"00",
													8585	=>X"00",
													8586	=>X"00",
													8587	=>X"00",
													8588	=>X"00",
													8589	=>X"00",
													8590	=>X"00",
													8591	=>X"00",
													8592	=>X"00",
													8593	=>X"00",
													8594	=>X"00",
													8595	=>X"00",
													8596	=>X"00",
													8597	=>X"00",
													8598	=>X"00",
													8599	=>X"00",
													8600	=>X"00",
													8601	=>X"00",
													8602	=>X"00",
													8603	=>X"00",
													8604	=>X"00",
													8605	=>X"00",
													8606	=>X"00",
													8607	=>X"00",
													8608	=>X"00",
													8609	=>X"00",
													8610	=>X"00",
													8611	=>X"00",
													8612	=>X"00",
													8613	=>X"00",
													8614	=>X"00",
													8615	=>X"00",
													8616	=>X"00",
													8617	=>X"00",
													8618	=>X"00",
													8619	=>X"00",
													8620	=>X"00",
													8621	=>X"00",
													8622	=>X"00",
													8623	=>X"00",
													8624	=>X"00",
													8625	=>X"00",
													8626	=>X"00",
													8627	=>X"00",
													8628	=>X"00",
													8629	=>X"00",
													8630	=>X"00",
													8631	=>X"00",
													8632	=>X"00",
													8633	=>X"00",
													8634	=>X"00",
													8635	=>X"00",
													8636	=>X"00",
													8637	=>X"00",
													8638	=>X"00",
													8639	=>X"00",
													8640	=>X"00",
													8641	=>X"00",
													8642	=>X"00",
													8643	=>X"00",
													8644	=>X"00",
													8645	=>X"00",
													8646	=>X"00",
													8647	=>X"00",
													8648	=>X"00",
													8649	=>X"00",
													8650	=>X"00",
													8651	=>X"00",
													8652	=>X"00",
													8653	=>X"00",
													8654	=>X"00",
													8655	=>X"00",
													8656	=>X"00",
													8657	=>X"00",
													8658	=>X"00",
													8659	=>X"00",
													8660	=>X"00",
													8661	=>X"00",
													8662	=>X"00",
													8663	=>X"00",
													8664	=>X"00",
													8665	=>X"00",
													8666	=>X"00",
													8667	=>X"00",
													8668	=>X"00",
													8669	=>X"00",
													8670	=>X"00",
													8671	=>X"00",
													8672	=>X"00",
													8673	=>X"00",
													8674	=>X"00",
													8675	=>X"00",
													8676	=>X"00",
													8677	=>X"00",
													8678	=>X"00",
													8679	=>X"00",
													8680	=>X"00",
													8681	=>X"00",
													8682	=>X"00",
													8683	=>X"00",
													8684	=>X"00",
													8685	=>X"00",
													8686	=>X"00",
													8687	=>X"00",
													8688	=>X"00",
													8689	=>X"00",
													8690	=>X"00",
													8691	=>X"00",
													8692	=>X"00",
													8693	=>X"00",
													8694	=>X"00",
													8695	=>X"00",
													8696	=>X"00",
													8697	=>X"00",
													8698	=>X"00",
													8699	=>X"00",
													8700	=>X"00",
													8701	=>X"00",
													8702	=>X"00",
													8703	=>X"00",
													8704	=>X"00",
													8705	=>X"00",
													8706	=>X"00",
													8707	=>X"00",
													8708	=>X"00",
													8709	=>X"00",
													8710	=>X"00",
													8711	=>X"00",
													8712	=>X"00",
													8713	=>X"00",
													8714	=>X"00",
													8715	=>X"00",
													8716	=>X"00",
													8717	=>X"00",
													8718	=>X"00",
													8719	=>X"00",
													8720	=>X"00",
													8721	=>X"00",
													8722	=>X"00",
													8723	=>X"00",
													8724	=>X"00",
													8725	=>X"00",
													8726	=>X"00",
													8727	=>X"00",
													8728	=>X"00",
													8729	=>X"00",
													8730	=>X"00",
													8731	=>X"00",
													8732	=>X"00",
													8733	=>X"00",
													8734	=>X"00",
													8735	=>X"00",
													8736	=>X"00",
													8737	=>X"00",
													8738	=>X"00",
													8739	=>X"00",
													8740	=>X"00",
													8741	=>X"00",
													8742	=>X"00",
													8743	=>X"00",
													8744	=>X"00",
													8745	=>X"00",
													8746	=>X"00",
													8747	=>X"00",
													8748	=>X"00",
													8749	=>X"00",
													8750	=>X"00",
													8751	=>X"00",
													8752	=>X"00",
													8753	=>X"00",
													8754	=>X"00",
													8755	=>X"00",
													8756	=>X"00",
													8757	=>X"00",
													8758	=>X"00",
													8759	=>X"00",
													8760	=>X"00",
													8761	=>X"00",
													8762	=>X"00",
													8763	=>X"00",
													8764	=>X"00",
													8765	=>X"00",
													8766	=>X"00",
													8767	=>X"00",
													8768	=>X"00",
													8769	=>X"00",
													8770	=>X"00",
													8771	=>X"00",
													8772	=>X"00",
													8773	=>X"00",
													8774	=>X"00",
													8775	=>X"00",
													8776	=>X"00",
													8777	=>X"00",
													8778	=>X"00",
													8779	=>X"00",
													8780	=>X"00",
													8781	=>X"00",
													8782	=>X"00",
													8783	=>X"00",
													8784	=>X"00",
													8785	=>X"00",
													8786	=>X"00",
													8787	=>X"00",
													8788	=>X"00",
													8789	=>X"00",
													8790	=>X"00",
													8791	=>X"00",
													8792	=>X"00",
													8793	=>X"00",
													8794	=>X"00",
													8795	=>X"00",
													8796	=>X"00",
													8797	=>X"00",
													8798	=>X"00",
													8799	=>X"00",
													8800	=>X"00",
													8801	=>X"00",
													8802	=>X"00",
													8803	=>X"00",
													8804	=>X"00",
													8805	=>X"00",
													8806	=>X"00",
													8807	=>X"00",
													8808	=>X"00",
													8809	=>X"00",
													8810	=>X"00",
													8811	=>X"00",
													8812	=>X"00",
													8813	=>X"00",
													8814	=>X"00",
													8815	=>X"00",
													8816	=>X"00",
													8817	=>X"00",
													8818	=>X"00",
													8819	=>X"00",
													8820	=>X"00",
													8821	=>X"00",
													8822	=>X"00",
													8823	=>X"00",
													8824	=>X"00",
													8825	=>X"00",
													8826	=>X"00",
													8827	=>X"00",
													8828	=>X"00",
													8829	=>X"00",
													8830	=>X"00",
													8831	=>X"00",
													8832	=>X"00",
													8833	=>X"00",
													8834	=>X"00",
													8835	=>X"00",
													8836	=>X"00",
													8837	=>X"00",
													8838	=>X"00",
													8839	=>X"00",
													8840	=>X"00",
													8841	=>X"00",
													8842	=>X"00",
													8843	=>X"00",
													8844	=>X"00",
													8845	=>X"00",
													8846	=>X"00",
													8847	=>X"00",
													8848	=>X"00",
													8849	=>X"00",
													8850	=>X"00",
													8851	=>X"00",
													8852	=>X"00",
													8853	=>X"00",
													8854	=>X"00",
													8855	=>X"00",
													8856	=>X"00",
													8857	=>X"00",
													8858	=>X"00",
													8859	=>X"00",
													8860	=>X"00",
													8861	=>X"00",
													8862	=>X"00",
													8863	=>X"00",
													8864	=>X"00",
													8865	=>X"00",
													8866	=>X"00",
													8867	=>X"00",
													8868	=>X"00",
													8869	=>X"00",
													8870	=>X"00",
													8871	=>X"00",
													8872	=>X"00",
													8873	=>X"00",
													8874	=>X"00",
													8875	=>X"00",
													8876	=>X"00",
													8877	=>X"00",
													8878	=>X"00",
													8879	=>X"00",
													8880	=>X"00",
													8881	=>X"00",
													8882	=>X"00",
													8883	=>X"00",
													8884	=>X"00",
													8885	=>X"00",
													8886	=>X"00",
													8887	=>X"00",
													8888	=>X"00",
													8889	=>X"00",
													8890	=>X"00",
													8891	=>X"00",
													8892	=>X"00",
													8893	=>X"00",
													8894	=>X"00",
													8895	=>X"00",
													8896	=>X"00",
													8897	=>X"00",
													8898	=>X"00",
													8899	=>X"00",
													8900	=>X"00",
													8901	=>X"00",
													8902	=>X"00",
													8903	=>X"00",
													8904	=>X"00",
													8905	=>X"00",
													8906	=>X"00",
													8907	=>X"00",
													8908	=>X"00",
													8909	=>X"00",
													8910	=>X"00",
													8911	=>X"00",
													8912	=>X"00",
													8913	=>X"00",
													8914	=>X"00",
													8915	=>X"00",
													8916	=>X"00",
													8917	=>X"00",
													8918	=>X"00",
													8919	=>X"00",
													8920	=>X"00",
													8921	=>X"00",
													8922	=>X"00",
													8923	=>X"00",
													8924	=>X"00",
													8925	=>X"00",
													8926	=>X"00",
													8927	=>X"00",
													8928	=>X"00",
													8929	=>X"00",
													8930	=>X"00",
													8931	=>X"00",
													8932	=>X"00",
													8933	=>X"00",
													8934	=>X"00",
													8935	=>X"00",
													8936	=>X"00",
													8937	=>X"00",
													8938	=>X"00",
													8939	=>X"00",
													8940	=>X"00",
													8941	=>X"00",
													8942	=>X"00",
													8943	=>X"00",
													8944	=>X"00",
													8945	=>X"00",
													8946	=>X"00",
													8947	=>X"00",
													8948	=>X"00",
													8949	=>X"00",
													8950	=>X"00",
													8951	=>X"00",
													8952	=>X"00",
													8953	=>X"00",
													8954	=>X"00",
													8955	=>X"00",
													8956	=>X"00",
													8957	=>X"00",
													8958	=>X"00",
													8959	=>X"00",
													8960	=>X"00",
													8961	=>X"00",
													8962	=>X"00",
													8963	=>X"00",
													8964	=>X"00",
													8965	=>X"00",
													8966	=>X"00",
													8967	=>X"00",
													8968	=>X"00",
													8969	=>X"00",
													8970	=>X"00",
													8971	=>X"00",
													8972	=>X"00",
													8973	=>X"00",
													8974	=>X"00",
													8975	=>X"00",
													8976	=>X"00",
													8977	=>X"00",
													8978	=>X"00",
													8979	=>X"00",
													8980	=>X"00",
													8981	=>X"00",
													8982	=>X"00",
													8983	=>X"00",
													8984	=>X"00",
													8985	=>X"00",
													8986	=>X"00",
													8987	=>X"00",
													8988	=>X"00",
													8989	=>X"00",
													8990	=>X"00",
													8991	=>X"00",
													8992	=>X"00",
													8993	=>X"00",
													8994	=>X"00",
													8995	=>X"00",
													8996	=>X"00",
													8997	=>X"00",
													8998	=>X"00",
													8999	=>X"00",
													9000	=>X"00",
													9001	=>X"00",
													9002	=>X"00",
													9003	=>X"00",
													9004	=>X"00",
													9005	=>X"00",
													9006	=>X"00",
													9007	=>X"00",
													9008	=>X"00",
													9009	=>X"00",
													9010	=>X"00",
													9011	=>X"00",
													9012	=>X"00",
													9013	=>X"00",
													9014	=>X"00",
													9015	=>X"00",
													9016	=>X"00",
													9017	=>X"00",
													9018	=>X"00",
													9019	=>X"00",
													9020	=>X"00",
													9021	=>X"00",
													9022	=>X"00",
													9023	=>X"00",
													9024	=>X"00",
													9025	=>X"00",
													9026	=>X"00",
													9027	=>X"00",
													9028	=>X"00",
													9029	=>X"00",
													9030	=>X"00",
													9031	=>X"00",
													9032	=>X"00",
													9033	=>X"00",
													9034	=>X"00",
													9035	=>X"00",
													9036	=>X"00",
													9037	=>X"00",
													9038	=>X"00",
													9039	=>X"00",
													9040	=>X"00",
													9041	=>X"00",
													9042	=>X"00",
													9043	=>X"00",
													9044	=>X"00",
													9045	=>X"00",
													9046	=>X"00",
													9047	=>X"00",
													9048	=>X"00",
													9049	=>X"00",
													9050	=>X"00",
													9051	=>X"00",
													9052	=>X"00",
													9053	=>X"00",
													9054	=>X"00",
													9055	=>X"00",
													9056	=>X"00",
													9057	=>X"00",
													9058	=>X"00",
													9059	=>X"00",
													9060	=>X"00",
													9061	=>X"00",
													9062	=>X"00",
													9063	=>X"00",
													9064	=>X"00",
													9065	=>X"00",
													9066	=>X"00",
													9067	=>X"00",
													9068	=>X"00",
													9069	=>X"00",
													9070	=>X"00",
													9071	=>X"00",
													9072	=>X"00",
													9073	=>X"00",
													9074	=>X"00",
													9075	=>X"00",
													9076	=>X"00",
													9077	=>X"00",
													9078	=>X"00",
													9079	=>X"00",
													9080	=>X"00",
													9081	=>X"00",
													9082	=>X"00",
													9083	=>X"00",
													9084	=>X"00",
													9085	=>X"00",
													9086	=>X"00",
													9087	=>X"00",
													9088	=>X"00",
													9089	=>X"00",
													9090	=>X"00",
													9091	=>X"00",
													9092	=>X"00",
													9093	=>X"00",
													9094	=>X"00",
													9095	=>X"00",
													9096	=>X"00",
													9097	=>X"00",
													9098	=>X"00",
													9099	=>X"00",
													9100	=>X"00",
													9101	=>X"00",
													9102	=>X"00",
													9103	=>X"00",
													9104	=>X"00",
													9105	=>X"00",
													9106	=>X"00",
													9107	=>X"00",
													9108	=>X"00",
													9109	=>X"00",
													9110	=>X"00",
													9111	=>X"00",
													9112	=>X"00",
													9113	=>X"00",
													9114	=>X"00",
													9115	=>X"00",
													9116	=>X"00",
													9117	=>X"00",
													9118	=>X"00",
													9119	=>X"00",
													9120	=>X"00",
													9121	=>X"00",
													9122	=>X"00",
													9123	=>X"00",
													9124	=>X"00",
													9125	=>X"00",
													9126	=>X"00",
													9127	=>X"00",
													9128	=>X"00",
													9129	=>X"00",
													9130	=>X"00",
													9131	=>X"00",
													9132	=>X"00",
													9133	=>X"00",
													9134	=>X"00",
													9135	=>X"00",
													9136	=>X"00",
													9137	=>X"00",
													9138	=>X"00",
													9139	=>X"00",
													9140	=>X"00",
													9141	=>X"00",
													9142	=>X"00",
													9143	=>X"00",
													9144	=>X"00",
													9145	=>X"00",
													9146	=>X"00",
													9147	=>X"00",
													9148	=>X"00",
													9149	=>X"00",
													9150	=>X"00",
													9151	=>X"00",
													9152	=>X"00",
													9153	=>X"00",
													9154	=>X"00",
													9155	=>X"00",
													9156	=>X"00",
													9157	=>X"00",
													9158	=>X"00",
													9159	=>X"00",
													9160	=>X"00",
													9161	=>X"00",
													9162	=>X"00",
													9163	=>X"00",
													9164	=>X"00",
													9165	=>X"00",
													9166	=>X"00",
													9167	=>X"00",
													9168	=>X"00",
													9169	=>X"00",
													9170	=>X"00",
													9171	=>X"00",
													9172	=>X"00",
													9173	=>X"00",
													9174	=>X"00",
													9175	=>X"00",
													9176	=>X"00",
													9177	=>X"00",
													9178	=>X"00",
													9179	=>X"00",
													9180	=>X"00",
													9181	=>X"00",
													9182	=>X"00",
													9183	=>X"00",
													9184	=>X"00",
													9185	=>X"00",
													9186	=>X"00",
													9187	=>X"00",
													9188	=>X"00",
													9189	=>X"00",
													9190	=>X"00",
													9191	=>X"00",
													9192	=>X"00",
													9193	=>X"00",
													9194	=>X"00",
													9195	=>X"00",
													9196	=>X"00",
													9197	=>X"00",
													9198	=>X"00",
													9199	=>X"00",
													9200	=>X"00",
													9201	=>X"00",
													9202	=>X"00",
													9203	=>X"00",
													9204	=>X"00",
													9205	=>X"00",
													9206	=>X"00",
													9207	=>X"00",
													9208	=>X"00",
													9209	=>X"00",
													9210	=>X"00",
													9211	=>X"00",
													9212	=>X"00",
													9213	=>X"00",
													9214	=>X"00",
													9215	=>X"00",
													9216	=>X"00",
													9217	=>X"00",
													9218	=>X"00",
													9219	=>X"00",
													9220	=>X"00",
													9221	=>X"00",
													9222	=>X"00",
													9223	=>X"00",
													9224	=>X"00",
													9225	=>X"00",
													9226	=>X"00",
													9227	=>X"00",
													9228	=>X"00",
													9229	=>X"00",
													9230	=>X"00",
													9231	=>X"00",
													9232	=>X"00",
													9233	=>X"00",
													9234	=>X"00",
													9235	=>X"00",
													9236	=>X"00",
													9237	=>X"00",
													9238	=>X"00",
													9239	=>X"00",
													9240	=>X"00",
													9241	=>X"00",
													9242	=>X"00",
													9243	=>X"00",
													9244	=>X"00",
													9245	=>X"00",
													9246	=>X"00",
													9247	=>X"00",
													9248	=>X"00",
													9249	=>X"00",
													9250	=>X"00",
													9251	=>X"00",
													9252	=>X"00",
													9253	=>X"00",
													9254	=>X"00",
													9255	=>X"00",
													9256	=>X"00",
													9257	=>X"00",
													9258	=>X"00",
													9259	=>X"00",
													9260	=>X"00",
													9261	=>X"00",
													9262	=>X"00",
													9263	=>X"00",
													9264	=>X"00",
													9265	=>X"00",
													9266	=>X"00",
													9267	=>X"00",
													9268	=>X"00",
													9269	=>X"00",
													9270	=>X"00",
													9271	=>X"00",
													9272	=>X"00",
													9273	=>X"00",
													9274	=>X"00",
													9275	=>X"00",
													9276	=>X"00",
													9277	=>X"00",
													9278	=>X"00",
													9279	=>X"00",
													9280	=>X"00",
													9281	=>X"00",
													9282	=>X"00",
													9283	=>X"00",
													9284	=>X"00",
													9285	=>X"00",
													9286	=>X"00",
													9287	=>X"00",
													9288	=>X"00",
													9289	=>X"00",
													9290	=>X"00",
													9291	=>X"00",
													9292	=>X"00",
													9293	=>X"00",
													9294	=>X"00",
													9295	=>X"00",
													9296	=>X"00",
													9297	=>X"00",
													9298	=>X"00",
													9299	=>X"00",
													9300	=>X"00",
													9301	=>X"00",
													9302	=>X"00",
													9303	=>X"00",
													9304	=>X"00",
													9305	=>X"00",
													9306	=>X"00",
													9307	=>X"00",
													9308	=>X"00",
													9309	=>X"00",
													9310	=>X"00",
													9311	=>X"00",
													9312	=>X"00",
													9313	=>X"00",
													9314	=>X"00",
													9315	=>X"00",
													9316	=>X"00",
													9317	=>X"00",
													9318	=>X"00",
													9319	=>X"00",
													9320	=>X"00",
													9321	=>X"00",
													9322	=>X"00",
													9323	=>X"00",
													9324	=>X"00",
													9325	=>X"00",
													9326	=>X"00",
													9327	=>X"00",
													9328	=>X"00",
													9329	=>X"00",
													9330	=>X"00",
													9331	=>X"00",
													9332	=>X"00",
													9333	=>X"00",
													9334	=>X"00",
													9335	=>X"00",
													9336	=>X"00",
													9337	=>X"00",
													9338	=>X"00",
													9339	=>X"00",
													9340	=>X"00",
													9341	=>X"00",
													9342	=>X"00",
													9343	=>X"00",
													9344	=>X"00",
													9345	=>X"00",
													9346	=>X"00",
													9347	=>X"00",
													9348	=>X"00",
													9349	=>X"00",
													9350	=>X"00",
													9351	=>X"00",
													9352	=>X"00",
													9353	=>X"00",
													9354	=>X"00",
													9355	=>X"00",
													9356	=>X"00",
													9357	=>X"00",
													9358	=>X"00",
													9359	=>X"00",
													9360	=>X"00",
													9361	=>X"00",
													9362	=>X"00",
													9363	=>X"00",
													9364	=>X"00",
													9365	=>X"00",
													9366	=>X"00",
													9367	=>X"00",
													9368	=>X"00",
													9369	=>X"00",
													9370	=>X"00",
													9371	=>X"00",
													9372	=>X"00",
													9373	=>X"00",
													9374	=>X"00",
													9375	=>X"00",
													9376	=>X"00",
													9377	=>X"00",
													9378	=>X"00",
													9379	=>X"00",
													9380	=>X"00",
													9381	=>X"00",
													9382	=>X"00",
													9383	=>X"00",
													9384	=>X"00",
													9385	=>X"00",
													9386	=>X"00",
													9387	=>X"00",
													9388	=>X"00",
													9389	=>X"00",
													9390	=>X"00",
													9391	=>X"00",
													9392	=>X"00",
													9393	=>X"00",
													9394	=>X"00",
													9395	=>X"00",
													9396	=>X"00",
													9397	=>X"00",
													9398	=>X"00",
													9399	=>X"00",
													9400	=>X"00",
													9401	=>X"00",
													9402	=>X"00",
													9403	=>X"00",
													9404	=>X"00",
													9405	=>X"00",
													9406	=>X"00",
													9407	=>X"00",
													9408	=>X"00",
													9409	=>X"00",
													9410	=>X"00",
													9411	=>X"00",
													9412	=>X"00",
													9413	=>X"00",
													9414	=>X"00",
													9415	=>X"00",
													9416	=>X"00",
													9417	=>X"00",
													9418	=>X"00",
													9419	=>X"00",
													9420	=>X"00",
													9421	=>X"00",
													9422	=>X"00",
													9423	=>X"00",
													9424	=>X"00",
													9425	=>X"00",
													9426	=>X"00",
													9427	=>X"00",
													9428	=>X"00",
													9429	=>X"00",
													9430	=>X"00",
													9431	=>X"00",
													9432	=>X"00",
													9433	=>X"00",
													9434	=>X"00",
													9435	=>X"00",
													9436	=>X"00",
													9437	=>X"00",
													9438	=>X"00",
													9439	=>X"00",
													9440	=>X"00",
													9441	=>X"00",
													9442	=>X"00",
													9443	=>X"00",
													9444	=>X"00",
													9445	=>X"00",
													9446	=>X"00",
													9447	=>X"00",
													9448	=>X"00",
													9449	=>X"00",
													9450	=>X"00",
													9451	=>X"00",
													9452	=>X"00",
													9453	=>X"00",
													9454	=>X"00",
													9455	=>X"00",
													9456	=>X"00",
													9457	=>X"00",
													9458	=>X"00",
													9459	=>X"00",
													9460	=>X"00",
													9461	=>X"00",
													9462	=>X"00",
													9463	=>X"00",
													9464	=>X"00",
													9465	=>X"00",
													9466	=>X"00",
													9467	=>X"00",
													9468	=>X"00",
													9469	=>X"00",
													9470	=>X"00",
													9471	=>X"00",
													9472	=>X"00",
													9473	=>X"00",
													9474	=>X"00",
													9475	=>X"00",
													9476	=>X"00",
													9477	=>X"00",
													9478	=>X"00",
													9479	=>X"00",
													9480	=>X"00",
													9481	=>X"00",
													9482	=>X"00",
													9483	=>X"00",
													9484	=>X"00",
													9485	=>X"00",
													9486	=>X"00",
													9487	=>X"00",
													9488	=>X"00",
													9489	=>X"00",
													9490	=>X"00",
													9491	=>X"00",
													9492	=>X"00",
													9493	=>X"00",
													9494	=>X"00",
													9495	=>X"00",
													9496	=>X"00",
													9497	=>X"00",
													9498	=>X"00",
													9499	=>X"00",
													9500	=>X"00",
													9501	=>X"00",
													9502	=>X"00",
													9503	=>X"00",
													9504	=>X"00",
													9505	=>X"00",
													9506	=>X"00",
													9507	=>X"00",
													9508	=>X"00",
													9509	=>X"00",
													9510	=>X"00",
													9511	=>X"00",
													9512	=>X"00",
													9513	=>X"00",
													9514	=>X"00",
													9515	=>X"00",
													9516	=>X"00",
													9517	=>X"00",
													9518	=>X"00",
													9519	=>X"00",
													9520	=>X"00",
													9521	=>X"00",
													9522	=>X"00",
													9523	=>X"00",
													9524	=>X"00",
													9525	=>X"00",
													9526	=>X"00",
													9527	=>X"00",
													9528	=>X"00",
													9529	=>X"00",
													9530	=>X"00",
													9531	=>X"00",
													9532	=>X"00",
													9533	=>X"00",
													9534	=>X"00",
													9535	=>X"00",
													9536	=>X"00",
													9537	=>X"00",
													9538	=>X"00",
													9539	=>X"00",
													9540	=>X"00",
													9541	=>X"00",
													9542	=>X"00",
													9543	=>X"00",
													9544	=>X"00",
													9545	=>X"00",
													9546	=>X"00",
													9547	=>X"00",
													9548	=>X"00",
													9549	=>X"00",
													9550	=>X"00",
													9551	=>X"00",
													9552	=>X"00",
													9553	=>X"00",
													9554	=>X"00",
													9555	=>X"00",
													9556	=>X"00",
													9557	=>X"00",
													9558	=>X"00",
													9559	=>X"00",
													9560	=>X"00",
													9561	=>X"00",
													9562	=>X"00",
													9563	=>X"00",
													9564	=>X"00",
													9565	=>X"00",
													9566	=>X"00",
													9567	=>X"00",
													9568	=>X"00",
													9569	=>X"00",
													9570	=>X"00",
													9571	=>X"00",
													9572	=>X"00",
													9573	=>X"00",
													9574	=>X"00",
													9575	=>X"00",
													9576	=>X"00",
													9577	=>X"00",
													9578	=>X"00",
													9579	=>X"00",
													9580	=>X"00",
													9581	=>X"00",
													9582	=>X"00",
													9583	=>X"00",
													9584	=>X"00",
													9585	=>X"00",
													9586	=>X"00",
													9587	=>X"00",
													9588	=>X"00",
													9589	=>X"00",
													9590	=>X"00",
													9591	=>X"00",
													9592	=>X"00",
													9593	=>X"00",
													9594	=>X"00",
													9595	=>X"00",
													9596	=>X"00",
													9597	=>X"00",
													9598	=>X"00",
													9599	=>X"00",
													9600	=>X"00",
													others=> X"00");	

									


signal sig_std_sys_set			:	std_logic := '0';
signal sig_std_scroll			:	std_logic := '0';
signal sig_std_hdot_scr			:	std_logic := '0';
signal sig_std_ovlay				:	std_logic := '0';

signal sig_std_disp_on			:	std_logic := '0';

signal sig_std_set_graph		:	std_logic := '0';
signal sig_std_clr_set_start	:	std_logic := '0';
signal sig_std_set_start		:	std_logic := '0';
signal sig_std_clr_disp			:	std_logic := '0';
signal sig_std_clr_graph		:	std_logic := '0';

signal sig_std_res				:	std_logic := '0';

signal sig_std_cgram_adr		:	std_logic := '0';
signal sig_std_draw_logo		: 	std_logic := '0';
signal sig_std_set_start_gr	:	std_logic := '0';



signal sig_std_init				: 	std_logic	:= '0';

signal sig_std8_start			: 	std_logic_vector(7 downto 0) := X"FF";
signal sig_test_data1			: 	std_logic_vector(255 downto 0);
signal sig_std_start				: 	std_logic							:='0';
signal sig_std_stop				: 	std_logic							:='0';
signal sig_std_strt				: 	std_logic							:='0';
signal sig_std_change_bit		:	std_logic							:='0';

signal sig_std_change_data		:	std_logic := '0';

signal sig_std_read_ok			: 	unsigned(11 downto 0);

signal sig_int_count				: 	integer	:=	0;
signal i 							: 	integer :=0;
signal sig_std_cmd 				: 	std_logic := '0';
signal sig_std_ready 			:	std_logic := '0';

signal sig_std_draw				:	std_logic	:=	'0';



signal sig_std_cnt 				:	integer := 0;
signal sig_int_numb_cnt			: 	integer := 0;


signal sig_std_lcd_mode				: std_logic	:=	'0';
signal var_int_cnt 				: integer := 0;


signal cur_arr : data (0 to 9600);
begin

out_std_oe_buf <= '1'	when (in_std_ena = '0') else
						'0';


WRK: process(in_std_ena,in_std_clk)

begin
	if (in_std_ena = '0') then
		sig_std_init	<=	'0';
		sig_std_res <= '0';
		var_int_cnt	<= 0;
		sig_std_sys_set <= '0';
		sig_std_scroll <= '0';
		sig_std_hdot_scr <= '0';
		sig_std_ovlay <= '0';
		sig_std_cgram_adr <= '0';
		sig_std_disp_on <= '0';
		sig_std_clr_disp <= '0';
		sig_std_clr_set_start <= '0';
		sig_std_draw <= '0';
		sig_std_set_start_gr <= '0';
		sig_std_set_start <= '0';
		sig_std_stop <= '0';
		
		
	elsif (in_std_clk'event and in_std_clk='1') then 
		if (sig_std_init= '0') then
			if (sig_std_res = '0') then
				if (var_int_cnt >= 0 and var_int_cnt <= 74) then
					var_int_cnt <= var_int_cnt + 1;
				elsif (var_int_cnt >= 75 and var_int_cnt <= 10149) then
					out_std_cs <= '0';
					out_std_wr <= '0';
					out_std_a <= '0';
					out_std7_data <= X"00";
					out_std_res <= '0';
					var_int_cnt <= var_int_cnt + 1;
				elsif (var_int_cnt >= 10150 and var_int_cnt <=20274) then
					out_std_res <= '1';
					out_std_cs <= '1';
					out_std_a <= '1';
					var_int_cnt <= var_int_cnt + 1;
				elsif (var_int_cnt = 20275) then
					var_int_cnt <= 0;
					sig_std_res <= '1';
				end if;
			elsif (sig_std_sys_set = '0') then
				write_cmd_data	(	out_std7_data,
									system_set(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(4),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_sys_set);

			elsif (sig_std_scroll = '0') then
				write_cmd_data	(	out_std7_data,
									scroll(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(6),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_scroll);
			elsif (sig_std_hdot_scr = '0') then
				write_cmd_data	(	out_std7_data,
									hdot_scr(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(1),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_hdot_scr);
			elsif (sig_std_ovlay = '0') then
				write_cmd_data	(	out_std7_data,
									ovlay(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(1),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_ovlay);
									
									
			elsif (sig_std_cgram_adr = '0') then
				write_cmd_data	(	out_std7_data,
									cgram_adr(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(2),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_cgram_adr);
									

			
			elsif (sig_std_disp_on = '0') then
					write_cmd_data	(	out_std7_data,
									disp_on(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(1),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_disp_on);
			
			elsif (sig_std_clr_disp = '0') then
				if (sig_std_clr_set_start = '0') then
					write_cmd_data	(	out_std7_data,
									set_start_clr(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(2),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_clr_set_start);
				else
					write_cmd_data	(	out_std7_data,
									clr_disp(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(8),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_clr_disp);
				end if;

			elsif (sig_std_draw = '0') then
				if (sig_std_set_start_gr = '0') then
					write_cmd_data	(	out_std7_data,
									set_start(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(2),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_set_start_gr);
				else
					write_cmd_data	(	out_std7_data,
									logo_elsiel(i),
									out_std_a,
									out_std_wr,
									out_std_cs,
									i,
									i_arr(7),
									sig_std_cnt,
									sig_std_cmd,
									sig_std_init);
				end if;
			end if;
			
		else
			if (sig_std_strt = '1') then
				if (sig_std_lcd_mode = '0') then
					if (sig_std_draw = '0') then
						if (sig_std_set_start = '0') then
							write_cmd_data	(	out_std7_data,
											set_start(i),
											out_std_a,
											out_std_wr,
											out_std_cs,
											i,
											i_arr(2),
											sig_std_cnt,
											sig_std_cmd,
											sig_std_set_start);
						else
							write_cmd_data	(	out_std7_data,
											logo_elsiel(i),
											out_std_a,
											out_std_wr,
											out_std_cs,
											i,
											i_arr(7),
											sig_std_cnt,
											sig_std_cmd,
											sig_std_stop);
						end if;
					end if;
				else
					if (sig_std_draw = '0') then
						if (sig_std_set_start = '0') then
							write_cmd_data	(	out_std7_data,
											set_start(i),
											out_std_a,
											out_std_wr,
											out_std_cs,
											i,
											i_arr(2),
											sig_std_cnt,
											sig_std_cmd,
											sig_std_set_start);
						else
							write_cmd_data	(	out_std7_data,
											cur_arr(i),
											out_std_a,
											out_std_wr,
											out_std_cs,
											i,
											i_arr(7),
											sig_std_cnt,
											sig_std_cmd,
											sig_std_stop);
						end if;
					end if;
				end if;
			else 
				sig_std_set_start <= '0';
				sig_std_draw <= '0';
				sig_std_stop <= '0';
				sig_std_lcd_mode <= in_std_lcd_mode;
			end if;
		end if;	
	end if;
end process; 
 
 
 



CNT_INT: process(in_std_ena,in_std_clk)
variable var_int_counter : integer range 0 to 25500000 := 0;
begin
		if (in_std_ena = '0') then
			var_int_counter := 0;
		elsif (in_std_clk'event and in_std_clk='1') then 
			if (sig_std_init= '1') then
				if (var_int_counter < 999999) then
					var_int_counter := var_int_counter + 1;
					sig_std_start <= '0';
				else 
					var_int_counter := 0;
					sig_std_start <= '1';
				end if;
			else
				var_int_counter := 0;
			end if;
		end if;
end process;



STROBE_start: process(in_std_ena,in_std_clk)

begin
		if (in_std_ena = '0') then
			
		elsif (in_std_clk'event and in_std_clk='1') then 
			if (sig_std_start = '1' and sig_std_start'last_value = '0') then
				sig_std_strt <= '1';
			elsif (sig_std_stop = '1' and sig_std_stop'last_value = '0') then
				sig_std_strt <= '0';
			end if;
		end if;
end process;


CUR_ARRAY: process(in_std_ena,in_std_clk)

begin
		if (in_std_ena = '0') then
			cur_arr (0) <= X"42";
		elsif (in_std_clk'event and in_std_clk='1') then 
			if (in_std_nwe = '0' and in_std_nwe'last_value = '1') then
				cur_arr((to_integer(unsigned(in_std16_adress)))) <= in_std8_data_in;
			else
			
			end if;
		end if;
end process;




CON: process(in_std_ena,in_std_clk)
variable var_int_counter : integer range 0 to 25500000 := 0;
begin
		if (in_std_ena = '0') then
			var_int_counter := 0;
		elsif (in_std_clk'event and in_std_clk='1') then 
				if (var_int_counter < 799999) then
					var_int_counter := var_int_counter + 1;
					out_std_str <= '0';
				else 
					var_int_counter := 0;
					out_std_str <= '1';
				end if;
		end if;
end process;



end LCD_ARCH;	
