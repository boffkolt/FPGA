-- terminal_qsys.vhd

-- Generated using ACDS version 16.1 203

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity terminal_qsys is
	port (
		base_addr_ddr_out_export                           : out   std_logic_vector(31 downto 0);                     --            base_addr_ddr_out.export
		clk_clk                                            : in    std_logic                      := '0';             --                          clk.clk
		control_out_export                                 : out   std_logic_vector(31 downto 0);                     --                  control_out.export
		hps_f2h_sdram0_data_address                        : in    std_logic_vector(26 downto 0)  := (others => '0'); --          hps_f2h_sdram0_data.address
		hps_f2h_sdram0_data_burstcount                     : in    std_logic_vector(7 downto 0)   := (others => '0'); --                             .burstcount
		hps_f2h_sdram0_data_waitrequest                    : out   std_logic;                                         --                             .waitrequest
		hps_f2h_sdram0_data_readdata                       : out   std_logic_vector(255 downto 0);                    --                             .readdata
		hps_f2h_sdram0_data_readdatavalid                  : out   std_logic;                                         --                             .readdatavalid
		hps_f2h_sdram0_data_read                           : in    std_logic                      := '0';             --                             .read
		hps_f2h_sdram0_data_writedata                      : in    std_logic_vector(255 downto 0) := (others => '0'); --                             .writedata
		hps_f2h_sdram0_data_byteenable                     : in    std_logic_vector(31 downto 0)  := (others => '0'); --                             .byteenable
		hps_f2h_sdram0_data_write                          : in    std_logic                      := '0';             --                             .write
		hps_f2h_stm_hw_events_stm_hwevents                 : in    std_logic_vector(27 downto 0)  := (others => '0'); --        hps_f2h_stm_hw_events.stm_hwevents
		hps_h2f_cold_reset_reset_n                         : out   std_logic;                                         --           hps_h2f_cold_reset.reset_n
		hps_h2f_warm_reset_handshake_h2f_pending_rst_req_n : out   std_logic;                                         -- hps_h2f_warm_reset_handshake.h2f_pending_rst_req_n
		hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n : in    std_logic                      := '0';             --                             .f2h_pending_rst_ack_n
		hps_hps_io_hps_io_emac1_inst_TX_CLK                : out   std_logic;                                         --                   hps_hps_io.hps_io_emac1_inst_TX_CLK
		hps_hps_io_hps_io_emac1_inst_TXD0                  : out   std_logic;                                         --                             .hps_io_emac1_inst_TXD0
		hps_hps_io_hps_io_emac1_inst_TXD1                  : out   std_logic;                                         --                             .hps_io_emac1_inst_TXD1
		hps_hps_io_hps_io_emac1_inst_TXD2                  : out   std_logic;                                         --                             .hps_io_emac1_inst_TXD2
		hps_hps_io_hps_io_emac1_inst_TXD3                  : out   std_logic;                                         --                             .hps_io_emac1_inst_TXD3
		hps_hps_io_hps_io_emac1_inst_RXD0                  : in    std_logic                      := '0';             --                             .hps_io_emac1_inst_RXD0
		hps_hps_io_hps_io_emac1_inst_MDIO                  : inout std_logic                      := '0';             --                             .hps_io_emac1_inst_MDIO
		hps_hps_io_hps_io_emac1_inst_MDC                   : out   std_logic;                                         --                             .hps_io_emac1_inst_MDC
		hps_hps_io_hps_io_emac1_inst_RX_CTL                : in    std_logic                      := '0';             --                             .hps_io_emac1_inst_RX_CTL
		hps_hps_io_hps_io_emac1_inst_TX_CTL                : out   std_logic;                                         --                             .hps_io_emac1_inst_TX_CTL
		hps_hps_io_hps_io_emac1_inst_RX_CLK                : in    std_logic                      := '0';             --                             .hps_io_emac1_inst_RX_CLK
		hps_hps_io_hps_io_emac1_inst_RXD1                  : in    std_logic                      := '0';             --                             .hps_io_emac1_inst_RXD1
		hps_hps_io_hps_io_emac1_inst_RXD2                  : in    std_logic                      := '0';             --                             .hps_io_emac1_inst_RXD2
		hps_hps_io_hps_io_emac1_inst_RXD3                  : in    std_logic                      := '0';             --                             .hps_io_emac1_inst_RXD3
		hps_hps_io_hps_io_sdio_inst_CMD                    : inout std_logic                      := '0';             --                             .hps_io_sdio_inst_CMD
		hps_hps_io_hps_io_sdio_inst_D0                     : inout std_logic                      := '0';             --                             .hps_io_sdio_inst_D0
		hps_hps_io_hps_io_sdio_inst_D1                     : inout std_logic                      := '0';             --                             .hps_io_sdio_inst_D1
		hps_hps_io_hps_io_sdio_inst_CLK                    : out   std_logic;                                         --                             .hps_io_sdio_inst_CLK
		hps_hps_io_hps_io_sdio_inst_D2                     : inout std_logic                      := '0';             --                             .hps_io_sdio_inst_D2
		hps_hps_io_hps_io_sdio_inst_D3                     : inout std_logic                      := '0';             --                             .hps_io_sdio_inst_D3
		hps_hps_io_hps_io_uart0_inst_RX                    : in    std_logic                      := '0';             --                             .hps_io_uart0_inst_RX
		hps_hps_io_hps_io_uart0_inst_TX                    : out   std_logic;                                         --                             .hps_io_uart0_inst_TX
		leds_out_export                                    : out   std_logic_vector(9 downto 0);                      --                     leds_out.export
		memory_mem_a                                       : out   std_logic_vector(14 downto 0);                     --                       memory.mem_a
		memory_mem_ba                                      : out   std_logic_vector(2 downto 0);                      --                             .mem_ba
		memory_mem_ck                                      : out   std_logic;                                         --                             .mem_ck
		memory_mem_ck_n                                    : out   std_logic;                                         --                             .mem_ck_n
		memory_mem_cke                                     : out   std_logic;                                         --                             .mem_cke
		memory_mem_cs_n                                    : out   std_logic;                                         --                             .mem_cs_n
		memory_mem_ras_n                                   : out   std_logic;                                         --                             .mem_ras_n
		memory_mem_cas_n                                   : out   std_logic;                                         --                             .mem_cas_n
		memory_mem_we_n                                    : out   std_logic;                                         --                             .mem_we_n
		memory_mem_reset_n                                 : out   std_logic;                                         --                             .mem_reset_n
		memory_mem_dq                                      : inout std_logic_vector(31 downto 0)  := (others => '0'); --                             .mem_dq
		memory_mem_dqs                                     : inout std_logic_vector(3 downto 0)   := (others => '0'); --                             .mem_dqs
		memory_mem_dqs_n                                   : inout std_logic_vector(3 downto 0)   := (others => '0'); --                             .mem_dqs_n
		memory_mem_odt                                     : out   std_logic;                                         --                             .mem_odt
		memory_mem_dm                                      : out   std_logic_vector(3 downto 0);                      --                             .mem_dm
		memory_oct_rzqin                                   : in    std_logic                      := '0';             --                             .oct_rzqin
		reset_reset_n                                      : in    std_logic                      := '0';             --                        reset.reset_n
		state_in_export                                    : in    std_logic_vector(31 downto 0)  := (others => '0'); --                     state_in.export
		switches_in_export                                 : in    std_logic_vector(9 downto 0)   := (others => '0')  --                  switches_in.export
	);
end entity terminal_qsys;

architecture rtl of terminal_qsys is
	component terminal_qsys_base_address_ddr is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component terminal_qsys_base_address_ddr;

	component terminal_qsys_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_cold_rst_n           : out   std_logic;                                         -- reset_n
			h2f_pending_rst_req_n    : out   std_logic;                                         -- h2f_pending_rst_req_n
			f2h_pending_rst_ack_n    : in    std_logic                      := 'X';             -- f2h_pending_rst_ack_n
			f2h_stm_hwevents         : in    std_logic_vector(27 downto 0)  := (others => 'X'); -- stm_hwevents
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			f2h_sdram0_clk           : in    std_logic                      := 'X';             -- clk
			f2h_sdram0_ADDRESS       : in    std_logic_vector(26 downto 0)  := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT    : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST   : out   std_logic;                                         -- waitrequest
			f2h_sdram0_READDATA      : out   std_logic_vector(255 downto 0);                    -- readdata
			f2h_sdram0_READDATAVALID : out   std_logic;                                         -- readdatavalid
			f2h_sdram0_READ          : in    std_logic                      := 'X';             -- read
			f2h_sdram0_WRITEDATA     : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE    : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE         : in    std_logic                      := 'X';             -- write
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_WSTRB                : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(31 downto 0);                     -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                          -- rready
		);
	end component terminal_qsys_hps;

	component terminal_qsys_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component terminal_qsys_leds;

	component terminal_qsys_rbf_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component terminal_qsys_rbf_id;

	component terminal_qsys_state is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component terminal_qsys_state;

	component terminal_qsys_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component terminal_qsys_switches;

	component terminal_qsys_mm_interconnect_0 is
		port (
			hps_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			rbf_id_reset_reset_bridge_in_reset_reset                          : in  std_logic                     := 'X';             -- reset
			base_address_ddr_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			base_address_ddr_s1_write                                         : out std_logic;                                        -- write
			base_address_ddr_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			base_address_ddr_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			base_address_ddr_s1_chipselect                                    : out std_logic;                                        -- chipselect
			control_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			control_s1_write                                                  : out std_logic;                                        -- write
			control_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			control_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			control_s1_chipselect                                             : out std_logic;                                        -- chipselect
			leds_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                                     : out std_logic;                                        -- write
			leds_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                                : out std_logic;                                        -- chipselect
			rbf_id_control_slave_address                                      : out std_logic_vector(0 downto 0);                     -- address
			rbf_id_control_slave_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			state_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			state_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			switches_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component terminal_qsys_mm_interconnect_0;

	component terminal_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component terminal_qsys_rst_controller;

	component terminal_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component terminal_qsys_rst_controller_001;

	signal hps_h2f_lw_axi_master_awburst                         : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_awburst
	signal hps_h2f_lw_axi_master_arlen                           : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_arlen
	signal hps_h2f_lw_axi_master_wstrb                           : std_logic_vector(3 downto 0);  -- hps:h2f_lw_WSTRB -> mm_interconnect_0:hps_h2f_lw_axi_master_wstrb
	signal hps_h2f_lw_axi_master_wready                          : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	signal hps_h2f_lw_axi_master_rid                             : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	signal hps_h2f_lw_axi_master_rready                          : std_logic;                     -- hps:h2f_lw_RREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_rready
	signal hps_h2f_lw_axi_master_awlen                           : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_awlen
	signal hps_h2f_lw_axi_master_wid                             : std_logic_vector(11 downto 0); -- hps:h2f_lw_WID -> mm_interconnect_0:hps_h2f_lw_axi_master_wid
	signal hps_h2f_lw_axi_master_arcache                         : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_arcache
	signal hps_h2f_lw_axi_master_wvalid                          : std_logic;                     -- hps:h2f_lw_WVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_wvalid
	signal hps_h2f_lw_axi_master_araddr                          : std_logic_vector(20 downto 0); -- hps:h2f_lw_ARADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_araddr
	signal hps_h2f_lw_axi_master_arprot                          : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_arprot
	signal hps_h2f_lw_axi_master_awprot                          : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_awprot
	signal hps_h2f_lw_axi_master_wdata                           : std_logic_vector(31 downto 0); -- hps:h2f_lw_WDATA -> mm_interconnect_0:hps_h2f_lw_axi_master_wdata
	signal hps_h2f_lw_axi_master_arvalid                         : std_logic;                     -- hps:h2f_lw_ARVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_arvalid
	signal hps_h2f_lw_axi_master_awcache                         : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_awcache
	signal hps_h2f_lw_axi_master_arid                            : std_logic_vector(11 downto 0); -- hps:h2f_lw_ARID -> mm_interconnect_0:hps_h2f_lw_axi_master_arid
	signal hps_h2f_lw_axi_master_arlock                          : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_arlock
	signal hps_h2f_lw_axi_master_awlock                          : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_awlock
	signal hps_h2f_lw_axi_master_awaddr                          : std_logic_vector(20 downto 0); -- hps:h2f_lw_AWADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_awaddr
	signal hps_h2f_lw_axi_master_bresp                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	signal hps_h2f_lw_axi_master_arready                         : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	signal hps_h2f_lw_axi_master_rdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	signal hps_h2f_lw_axi_master_awready                         : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	signal hps_h2f_lw_axi_master_arburst                         : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_arburst
	signal hps_h2f_lw_axi_master_arsize                          : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_arsize
	signal hps_h2f_lw_axi_master_bready                          : std_logic;                     -- hps:h2f_lw_BREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_bready
	signal hps_h2f_lw_axi_master_rlast                           : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	signal hps_h2f_lw_axi_master_wlast                           : std_logic;                     -- hps:h2f_lw_WLAST -> mm_interconnect_0:hps_h2f_lw_axi_master_wlast
	signal hps_h2f_lw_axi_master_rresp                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	signal hps_h2f_lw_axi_master_awid                            : std_logic_vector(11 downto 0); -- hps:h2f_lw_AWID -> mm_interconnect_0:hps_h2f_lw_axi_master_awid
	signal hps_h2f_lw_axi_master_bid                             : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	signal hps_h2f_lw_axi_master_bvalid                          : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	signal hps_h2f_lw_axi_master_awsize                          : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_awsize
	signal hps_h2f_lw_axi_master_awvalid                         : std_logic;                     -- hps:h2f_lw_AWVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_awvalid
	signal hps_h2f_lw_axi_master_rvalid                          : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	signal mm_interconnect_0_rbf_id_control_slave_readdata       : std_logic_vector(31 downto 0); -- rbf_id:readdata -> mm_interconnect_0:rbf_id_control_slave_readdata
	signal mm_interconnect_0_rbf_id_control_slave_address        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:rbf_id_control_slave_address -> rbf_id:address
	signal mm_interconnect_0_state_s1_readdata                   : std_logic_vector(31 downto 0); -- state:readdata -> mm_interconnect_0:state_s1_readdata
	signal mm_interconnect_0_state_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:state_s1_address -> state:address
	signal mm_interconnect_0_control_s1_chipselect               : std_logic;                     -- mm_interconnect_0:control_s1_chipselect -> control:chipselect
	signal mm_interconnect_0_control_s1_readdata                 : std_logic_vector(31 downto 0); -- control:readdata -> mm_interconnect_0:control_s1_readdata
	signal mm_interconnect_0_control_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:control_s1_address -> control:address
	signal mm_interconnect_0_control_s1_write                    : std_logic;                     -- mm_interconnect_0:control_s1_write -> mm_interconnect_0_control_s1_write:in
	signal mm_interconnect_0_control_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:control_s1_writedata -> control:writedata
	signal mm_interconnect_0_base_address_ddr_s1_chipselect      : std_logic;                     -- mm_interconnect_0:base_address_ddr_s1_chipselect -> base_address_ddr:chipselect
	signal mm_interconnect_0_base_address_ddr_s1_readdata        : std_logic_vector(31 downto 0); -- base_address_ddr:readdata -> mm_interconnect_0:base_address_ddr_s1_readdata
	signal mm_interconnect_0_base_address_ddr_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:base_address_ddr_s1_address -> base_address_ddr:address
	signal mm_interconnect_0_base_address_ddr_s1_write           : std_logic;                     -- mm_interconnect_0:base_address_ddr_s1_write -> mm_interconnect_0_base_address_ddr_s1_write:in
	signal mm_interconnect_0_base_address_ddr_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:base_address_ddr_s1_writedata -> base_address_ddr:writedata
	signal mm_interconnect_0_leds_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                    : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                       : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_switches_s1_readdata                : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal rst_controller_reset_out_reset                        : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:rbf_id_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal hps_h2f_reset_reset                                   : std_logic;                     -- hps:h2f_rst_n -> hps_h2f_reset_reset:in
	signal rst_controller_001_reset_out_reset                    : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_0:hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal reset_reset_n_ports_inv                               : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_control_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_0_control_s1_write:inv -> control:write_n
	signal mm_interconnect_0_base_address_ddr_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_base_address_ddr_s1_write:inv -> base_address_ddr:write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal rst_controller_reset_out_reset_ports_inv              : std_logic;                     -- rst_controller_reset_out_reset:inv -> [base_address_ddr:reset_n, control:reset_n, leds:reset_n, rbf_id:reset_n, state:reset_n, switches:reset_n]
	signal hps_h2f_reset_reset_ports_inv                         : std_logic;                     -- hps_h2f_reset_reset:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in0]

begin

	base_address_ddr : component terminal_qsys_base_address_ddr
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_base_address_ddr_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_base_address_ddr_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_base_address_ddr_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_base_address_ddr_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_base_address_ddr_s1_readdata,        --                    .readdata
			out_port   => base_addr_ddr_out_export                               -- external_connection.export
		);

	control : component terminal_qsys_base_address_ddr
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_control_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_control_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_control_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_control_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_control_s1_readdata,        --                    .readdata
			out_port   => control_out_export                            -- external_connection.export
		);

	hps : component terminal_qsys_hps
		generic map (
			F2S_Width => 1,
			S2F_Width => 1
		)
		port map (
			h2f_cold_rst_n           => hps_h2f_cold_reset_reset_n,                         --           h2f_cold_reset.reset_n
			h2f_pending_rst_req_n    => hps_h2f_warm_reset_handshake_h2f_pending_rst_req_n, -- h2f_warm_reset_handshake.h2f_pending_rst_req_n
			f2h_pending_rst_ack_n    => hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n, --                         .f2h_pending_rst_ack_n
			f2h_stm_hwevents         => hps_f2h_stm_hw_events_stm_hwevents,                 --        f2h_stm_hw_events.stm_hwevents
			mem_a                    => memory_mem_a,                                       --                   memory.mem_a
			mem_ba                   => memory_mem_ba,                                      --                         .mem_ba
			mem_ck                   => memory_mem_ck,                                      --                         .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                                    --                         .mem_ck_n
			mem_cke                  => memory_mem_cke,                                     --                         .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                                    --                         .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                                   --                         .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                                   --                         .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                                    --                         .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                                 --                         .mem_reset_n
			mem_dq                   => memory_mem_dq,                                      --                         .mem_dq
			mem_dqs                  => memory_mem_dqs,                                     --                         .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                                   --                         .mem_dqs_n
			mem_odt                  => memory_mem_odt,                                     --                         .mem_odt
			mem_dm                   => memory_mem_dm,                                      --                         .mem_dm
			oct_rzqin                => memory_oct_rzqin,                                   --                         .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_hps_io_hps_io_emac1_inst_TX_CLK,                --                   hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_hps_io_hps_io_emac1_inst_TXD0,                  --                         .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_hps_io_hps_io_emac1_inst_TXD1,                  --                         .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_hps_io_hps_io_emac1_inst_TXD2,                  --                         .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_hps_io_hps_io_emac1_inst_TXD3,                  --                         .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_hps_io_hps_io_emac1_inst_RXD0,                  --                         .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_hps_io_hps_io_emac1_inst_MDIO,                  --                         .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_hps_io_hps_io_emac1_inst_MDC,                   --                         .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_hps_io_hps_io_emac1_inst_RX_CTL,                --                         .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_hps_io_hps_io_emac1_inst_TX_CTL,                --                         .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_hps_io_hps_io_emac1_inst_RX_CLK,                --                         .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_hps_io_hps_io_emac1_inst_RXD1,                  --                         .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_hps_io_hps_io_emac1_inst_RXD2,                  --                         .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_hps_io_hps_io_emac1_inst_RXD3,                  --                         .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_hps_io_hps_io_sdio_inst_CMD,                    --                         .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_hps_io_hps_io_sdio_inst_D0,                     --                         .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_hps_io_hps_io_sdio_inst_D1,                     --                         .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_hps_io_hps_io_sdio_inst_CLK,                    --                         .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_hps_io_hps_io_sdio_inst_D2,                     --                         .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_hps_io_hps_io_sdio_inst_D3,                     --                         .hps_io_sdio_inst_D3
			hps_io_uart0_inst_RX     => hps_hps_io_hps_io_uart0_inst_RX,                    --                         .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_hps_io_hps_io_uart0_inst_TX,                    --                         .hps_io_uart0_inst_TX
			h2f_rst_n                => hps_h2f_reset_reset,                                --                h2f_reset.reset_n
			f2h_sdram0_clk           => clk_clk,                                            --         f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS       => hps_f2h_sdram0_data_address,                        --          f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT    => hps_f2h_sdram0_data_burstcount,                     --                         .burstcount
			f2h_sdram0_WAITREQUEST   => hps_f2h_sdram0_data_waitrequest,                    --                         .waitrequest
			f2h_sdram0_READDATA      => hps_f2h_sdram0_data_readdata,                       --                         .readdata
			f2h_sdram0_READDATAVALID => hps_f2h_sdram0_data_readdatavalid,                  --                         .readdatavalid
			f2h_sdram0_READ          => hps_f2h_sdram0_data_read,                           --                         .read
			f2h_sdram0_WRITEDATA     => hps_f2h_sdram0_data_writedata,                      --                         .writedata
			f2h_sdram0_BYTEENABLE    => hps_f2h_sdram0_data_byteenable,                     --                         .byteenable
			f2h_sdram0_WRITE         => hps_f2h_sdram0_data_write,                          --                         .write
			h2f_axi_clk              => clk_clk,                                            --            h2f_axi_clock.clk
			h2f_AWID                 => open,                                               --           h2f_axi_master.awid
			h2f_AWADDR               => open,                                               --                         .awaddr
			h2f_AWLEN                => open,                                               --                         .awlen
			h2f_AWSIZE               => open,                                               --                         .awsize
			h2f_AWBURST              => open,                                               --                         .awburst
			h2f_AWLOCK               => open,                                               --                         .awlock
			h2f_AWCACHE              => open,                                               --                         .awcache
			h2f_AWPROT               => open,                                               --                         .awprot
			h2f_AWVALID              => open,                                               --                         .awvalid
			h2f_AWREADY              => open,                                               --                         .awready
			h2f_WID                  => open,                                               --                         .wid
			h2f_WDATA                => open,                                               --                         .wdata
			h2f_WSTRB                => open,                                               --                         .wstrb
			h2f_WLAST                => open,                                               --                         .wlast
			h2f_WVALID               => open,                                               --                         .wvalid
			h2f_WREADY               => open,                                               --                         .wready
			h2f_BID                  => open,                                               --                         .bid
			h2f_BRESP                => open,                                               --                         .bresp
			h2f_BVALID               => open,                                               --                         .bvalid
			h2f_BREADY               => open,                                               --                         .bready
			h2f_ARID                 => open,                                               --                         .arid
			h2f_ARADDR               => open,                                               --                         .araddr
			h2f_ARLEN                => open,                                               --                         .arlen
			h2f_ARSIZE               => open,                                               --                         .arsize
			h2f_ARBURST              => open,                                               --                         .arburst
			h2f_ARLOCK               => open,                                               --                         .arlock
			h2f_ARCACHE              => open,                                               --                         .arcache
			h2f_ARPROT               => open,                                               --                         .arprot
			h2f_ARVALID              => open,                                               --                         .arvalid
			h2f_ARREADY              => open,                                               --                         .arready
			h2f_RID                  => open,                                               --                         .rid
			h2f_RDATA                => open,                                               --                         .rdata
			h2f_RRESP                => open,                                               --                         .rresp
			h2f_RLAST                => open,                                               --                         .rlast
			h2f_RVALID               => open,                                               --                         .rvalid
			h2f_RREADY               => open,                                               --                         .rready
			f2h_axi_clk              => clk_clk,                                            --            f2h_axi_clock.clk
			f2h_AWID                 => open,                                               --            f2h_axi_slave.awid
			f2h_AWADDR               => open,                                               --                         .awaddr
			f2h_AWLEN                => open,                                               --                         .awlen
			f2h_AWSIZE               => open,                                               --                         .awsize
			f2h_AWBURST              => open,                                               --                         .awburst
			f2h_AWLOCK               => open,                                               --                         .awlock
			f2h_AWCACHE              => open,                                               --                         .awcache
			f2h_AWPROT               => open,                                               --                         .awprot
			f2h_AWVALID              => open,                                               --                         .awvalid
			f2h_AWREADY              => open,                                               --                         .awready
			f2h_AWUSER               => open,                                               --                         .awuser
			f2h_WID                  => open,                                               --                         .wid
			f2h_WDATA                => open,                                               --                         .wdata
			f2h_WSTRB                => open,                                               --                         .wstrb
			f2h_WLAST                => open,                                               --                         .wlast
			f2h_WVALID               => open,                                               --                         .wvalid
			f2h_WREADY               => open,                                               --                         .wready
			f2h_BID                  => open,                                               --                         .bid
			f2h_BRESP                => open,                                               --                         .bresp
			f2h_BVALID               => open,                                               --                         .bvalid
			f2h_BREADY               => open,                                               --                         .bready
			f2h_ARID                 => open,                                               --                         .arid
			f2h_ARADDR               => open,                                               --                         .araddr
			f2h_ARLEN                => open,                                               --                         .arlen
			f2h_ARSIZE               => open,                                               --                         .arsize
			f2h_ARBURST              => open,                                               --                         .arburst
			f2h_ARLOCK               => open,                                               --                         .arlock
			f2h_ARCACHE              => open,                                               --                         .arcache
			f2h_ARPROT               => open,                                               --                         .arprot
			f2h_ARVALID              => open,                                               --                         .arvalid
			f2h_ARREADY              => open,                                               --                         .arready
			f2h_ARUSER               => open,                                               --                         .aruser
			f2h_RID                  => open,                                               --                         .rid
			f2h_RDATA                => open,                                               --                         .rdata
			f2h_RRESP                => open,                                               --                         .rresp
			f2h_RLAST                => open,                                               --                         .rlast
			f2h_RVALID               => open,                                               --                         .rvalid
			f2h_RREADY               => open,                                               --                         .rready
			h2f_lw_axi_clk           => clk_clk,                                            --         h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_h2f_lw_axi_master_awid,                         --        h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_h2f_lw_axi_master_awaddr,                       --                         .awaddr
			h2f_lw_AWLEN             => hps_h2f_lw_axi_master_awlen,                        --                         .awlen
			h2f_lw_AWSIZE            => hps_h2f_lw_axi_master_awsize,                       --                         .awsize
			h2f_lw_AWBURST           => hps_h2f_lw_axi_master_awburst,                      --                         .awburst
			h2f_lw_AWLOCK            => hps_h2f_lw_axi_master_awlock,                       --                         .awlock
			h2f_lw_AWCACHE           => hps_h2f_lw_axi_master_awcache,                      --                         .awcache
			h2f_lw_AWPROT            => hps_h2f_lw_axi_master_awprot,                       --                         .awprot
			h2f_lw_AWVALID           => hps_h2f_lw_axi_master_awvalid,                      --                         .awvalid
			h2f_lw_AWREADY           => hps_h2f_lw_axi_master_awready,                      --                         .awready
			h2f_lw_WID               => hps_h2f_lw_axi_master_wid,                          --                         .wid
			h2f_lw_WDATA             => hps_h2f_lw_axi_master_wdata,                        --                         .wdata
			h2f_lw_WSTRB             => hps_h2f_lw_axi_master_wstrb,                        --                         .wstrb
			h2f_lw_WLAST             => hps_h2f_lw_axi_master_wlast,                        --                         .wlast
			h2f_lw_WVALID            => hps_h2f_lw_axi_master_wvalid,                       --                         .wvalid
			h2f_lw_WREADY            => hps_h2f_lw_axi_master_wready,                       --                         .wready
			h2f_lw_BID               => hps_h2f_lw_axi_master_bid,                          --                         .bid
			h2f_lw_BRESP             => hps_h2f_lw_axi_master_bresp,                        --                         .bresp
			h2f_lw_BVALID            => hps_h2f_lw_axi_master_bvalid,                       --                         .bvalid
			h2f_lw_BREADY            => hps_h2f_lw_axi_master_bready,                       --                         .bready
			h2f_lw_ARID              => hps_h2f_lw_axi_master_arid,                         --                         .arid
			h2f_lw_ARADDR            => hps_h2f_lw_axi_master_araddr,                       --                         .araddr
			h2f_lw_ARLEN             => hps_h2f_lw_axi_master_arlen,                        --                         .arlen
			h2f_lw_ARSIZE            => hps_h2f_lw_axi_master_arsize,                       --                         .arsize
			h2f_lw_ARBURST           => hps_h2f_lw_axi_master_arburst,                      --                         .arburst
			h2f_lw_ARLOCK            => hps_h2f_lw_axi_master_arlock,                       --                         .arlock
			h2f_lw_ARCACHE           => hps_h2f_lw_axi_master_arcache,                      --                         .arcache
			h2f_lw_ARPROT            => hps_h2f_lw_axi_master_arprot,                       --                         .arprot
			h2f_lw_ARVALID           => hps_h2f_lw_axi_master_arvalid,                      --                         .arvalid
			h2f_lw_ARREADY           => hps_h2f_lw_axi_master_arready,                      --                         .arready
			h2f_lw_RID               => hps_h2f_lw_axi_master_rid,                          --                         .rid
			h2f_lw_RDATA             => hps_h2f_lw_axi_master_rdata,                        --                         .rdata
			h2f_lw_RRESP             => hps_h2f_lw_axi_master_rresp,                        --                         .rresp
			h2f_lw_RLAST             => hps_h2f_lw_axi_master_rlast,                        --                         .rlast
			h2f_lw_RVALID            => hps_h2f_lw_axi_master_rvalid,                       --                         .rvalid
			h2f_lw_RREADY            => hps_h2f_lw_axi_master_rready                        --                         .rready
		);

	leds : component terminal_qsys_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_out_export                            -- external_connection.export
		);

	rbf_id : component terminal_qsys_rbf_id
		port map (
			clock    => clk_clk,                                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_rbf_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_rbf_id_control_slave_address(0)  --              .address
		);

	state : component terminal_qsys_state
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_state_s1_address,       --                  s1.address
			readdata => mm_interconnect_0_state_s1_readdata,      --                    .readdata
			in_port  => state_in_export                           -- external_connection.export
		);

	switches : component terminal_qsys_switches
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,   --                    .readdata
			in_port  => switches_in_export                        -- external_connection.export
		);

	mm_interconnect_0 : component terminal_qsys_mm_interconnect_0
		port map (
			hps_h2f_lw_axi_master_awid                                        => hps_h2f_lw_axi_master_awid,                       --                                       hps_h2f_lw_axi_master.awid
			hps_h2f_lw_axi_master_awaddr                                      => hps_h2f_lw_axi_master_awaddr,                     --                                                            .awaddr
			hps_h2f_lw_axi_master_awlen                                       => hps_h2f_lw_axi_master_awlen,                      --                                                            .awlen
			hps_h2f_lw_axi_master_awsize                                      => hps_h2f_lw_axi_master_awsize,                     --                                                            .awsize
			hps_h2f_lw_axi_master_awburst                                     => hps_h2f_lw_axi_master_awburst,                    --                                                            .awburst
			hps_h2f_lw_axi_master_awlock                                      => hps_h2f_lw_axi_master_awlock,                     --                                                            .awlock
			hps_h2f_lw_axi_master_awcache                                     => hps_h2f_lw_axi_master_awcache,                    --                                                            .awcache
			hps_h2f_lw_axi_master_awprot                                      => hps_h2f_lw_axi_master_awprot,                     --                                                            .awprot
			hps_h2f_lw_axi_master_awvalid                                     => hps_h2f_lw_axi_master_awvalid,                    --                                                            .awvalid
			hps_h2f_lw_axi_master_awready                                     => hps_h2f_lw_axi_master_awready,                    --                                                            .awready
			hps_h2f_lw_axi_master_wid                                         => hps_h2f_lw_axi_master_wid,                        --                                                            .wid
			hps_h2f_lw_axi_master_wdata                                       => hps_h2f_lw_axi_master_wdata,                      --                                                            .wdata
			hps_h2f_lw_axi_master_wstrb                                       => hps_h2f_lw_axi_master_wstrb,                      --                                                            .wstrb
			hps_h2f_lw_axi_master_wlast                                       => hps_h2f_lw_axi_master_wlast,                      --                                                            .wlast
			hps_h2f_lw_axi_master_wvalid                                      => hps_h2f_lw_axi_master_wvalid,                     --                                                            .wvalid
			hps_h2f_lw_axi_master_wready                                      => hps_h2f_lw_axi_master_wready,                     --                                                            .wready
			hps_h2f_lw_axi_master_bid                                         => hps_h2f_lw_axi_master_bid,                        --                                                            .bid
			hps_h2f_lw_axi_master_bresp                                       => hps_h2f_lw_axi_master_bresp,                      --                                                            .bresp
			hps_h2f_lw_axi_master_bvalid                                      => hps_h2f_lw_axi_master_bvalid,                     --                                                            .bvalid
			hps_h2f_lw_axi_master_bready                                      => hps_h2f_lw_axi_master_bready,                     --                                                            .bready
			hps_h2f_lw_axi_master_arid                                        => hps_h2f_lw_axi_master_arid,                       --                                                            .arid
			hps_h2f_lw_axi_master_araddr                                      => hps_h2f_lw_axi_master_araddr,                     --                                                            .araddr
			hps_h2f_lw_axi_master_arlen                                       => hps_h2f_lw_axi_master_arlen,                      --                                                            .arlen
			hps_h2f_lw_axi_master_arsize                                      => hps_h2f_lw_axi_master_arsize,                     --                                                            .arsize
			hps_h2f_lw_axi_master_arburst                                     => hps_h2f_lw_axi_master_arburst,                    --                                                            .arburst
			hps_h2f_lw_axi_master_arlock                                      => hps_h2f_lw_axi_master_arlock,                     --                                                            .arlock
			hps_h2f_lw_axi_master_arcache                                     => hps_h2f_lw_axi_master_arcache,                    --                                                            .arcache
			hps_h2f_lw_axi_master_arprot                                      => hps_h2f_lw_axi_master_arprot,                     --                                                            .arprot
			hps_h2f_lw_axi_master_arvalid                                     => hps_h2f_lw_axi_master_arvalid,                    --                                                            .arvalid
			hps_h2f_lw_axi_master_arready                                     => hps_h2f_lw_axi_master_arready,                    --                                                            .arready
			hps_h2f_lw_axi_master_rid                                         => hps_h2f_lw_axi_master_rid,                        --                                                            .rid
			hps_h2f_lw_axi_master_rdata                                       => hps_h2f_lw_axi_master_rdata,                      --                                                            .rdata
			hps_h2f_lw_axi_master_rresp                                       => hps_h2f_lw_axi_master_rresp,                      --                                                            .rresp
			hps_h2f_lw_axi_master_rlast                                       => hps_h2f_lw_axi_master_rlast,                      --                                                            .rlast
			hps_h2f_lw_axi_master_rvalid                                      => hps_h2f_lw_axi_master_rvalid,                     --                                                            .rvalid
			hps_h2f_lw_axi_master_rready                                      => hps_h2f_lw_axi_master_rready,                     --                                                            .rready
			clk_clk_clk                                                       => clk_clk,                                          --                                                     clk_clk.clk
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,               -- hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			rbf_id_reset_reset_bridge_in_reset_reset                          => rst_controller_reset_out_reset,                   --                          rbf_id_reset_reset_bridge_in_reset.reset
			base_address_ddr_s1_address                                       => mm_interconnect_0_base_address_ddr_s1_address,    --                                         base_address_ddr_s1.address
			base_address_ddr_s1_write                                         => mm_interconnect_0_base_address_ddr_s1_write,      --                                                            .write
			base_address_ddr_s1_readdata                                      => mm_interconnect_0_base_address_ddr_s1_readdata,   --                                                            .readdata
			base_address_ddr_s1_writedata                                     => mm_interconnect_0_base_address_ddr_s1_writedata,  --                                                            .writedata
			base_address_ddr_s1_chipselect                                    => mm_interconnect_0_base_address_ddr_s1_chipselect, --                                                            .chipselect
			control_s1_address                                                => mm_interconnect_0_control_s1_address,             --                                                  control_s1.address
			control_s1_write                                                  => mm_interconnect_0_control_s1_write,               --                                                            .write
			control_s1_readdata                                               => mm_interconnect_0_control_s1_readdata,            --                                                            .readdata
			control_s1_writedata                                              => mm_interconnect_0_control_s1_writedata,           --                                                            .writedata
			control_s1_chipselect                                             => mm_interconnect_0_control_s1_chipselect,          --                                                            .chipselect
			leds_s1_address                                                   => mm_interconnect_0_leds_s1_address,                --                                                     leds_s1.address
			leds_s1_write                                                     => mm_interconnect_0_leds_s1_write,                  --                                                            .write
			leds_s1_readdata                                                  => mm_interconnect_0_leds_s1_readdata,               --                                                            .readdata
			leds_s1_writedata                                                 => mm_interconnect_0_leds_s1_writedata,              --                                                            .writedata
			leds_s1_chipselect                                                => mm_interconnect_0_leds_s1_chipselect,             --                                                            .chipselect
			rbf_id_control_slave_address                                      => mm_interconnect_0_rbf_id_control_slave_address,   --                                        rbf_id_control_slave.address
			rbf_id_control_slave_readdata                                     => mm_interconnect_0_rbf_id_control_slave_readdata,  --                                                            .readdata
			state_s1_address                                                  => mm_interconnect_0_state_s1_address,               --                                                    state_s1.address
			state_s1_readdata                                                 => mm_interconnect_0_state_s1_readdata,              --                                                            .readdata
			switches_s1_address                                               => mm_interconnect_0_switches_s1_address,            --                                                 switches_s1.address
			switches_s1_readdata                                              => mm_interconnect_0_switches_s1_readdata            --                                                            .readdata
		);

	rst_controller : component terminal_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			reset_in1      => hps_h2f_reset_reset_ports_inv,  -- reset_in1.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component terminal_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_h2f_reset_reset_ports_inv,      -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_control_s1_write_ports_inv <= not mm_interconnect_0_control_s1_write;

	mm_interconnect_0_base_address_ddr_s1_write_ports_inv <= not mm_interconnect_0_base_address_ddr_s1_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_h2f_reset_reset_ports_inv <= not hps_h2f_reset_reset;

end architecture rtl; -- of terminal_qsys
