// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 16.1.2 Build 203 01/18/2017 SJ Lite Edition"

// DATE "06/07/2017 17:37:52"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module terminal_qsys (
	base_addr_ddr_out_export,
	clk_clk,
	control_out_export,
	hps_f2h_sdram0_data_address,
	hps_f2h_sdram0_data_burstcount,
	hps_f2h_sdram0_data_waitrequest,
	hps_f2h_sdram0_data_readdata,
	hps_f2h_sdram0_data_readdatavalid,
	hps_f2h_sdram0_data_read,
	hps_f2h_sdram0_data_writedata,
	hps_f2h_sdram0_data_byteenable,
	hps_f2h_sdram0_data_write,
	hps_f2h_stm_hw_events_stm_hwevents,
	hps_h2f_cold_reset_reset_n,
	hps_h2f_warm_reset_handshake_h2f_pending_rst_req_n,
	hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n,
	hps_hps_io_hps_io_emac1_inst_TX_CLK,
	hps_hps_io_hps_io_emac1_inst_TXD0,
	hps_hps_io_hps_io_emac1_inst_TXD1,
	hps_hps_io_hps_io_emac1_inst_TXD2,
	hps_hps_io_hps_io_emac1_inst_TXD3,
	hps_hps_io_hps_io_emac1_inst_RXD0,
	hps_hps_io_hps_io_emac1_inst_MDIO,
	hps_hps_io_hps_io_emac1_inst_MDC,
	hps_hps_io_hps_io_emac1_inst_RX_CTL,
	hps_hps_io_hps_io_emac1_inst_TX_CTL,
	hps_hps_io_hps_io_emac1_inst_RX_CLK,
	hps_hps_io_hps_io_emac1_inst_RXD1,
	hps_hps_io_hps_io_emac1_inst_RXD2,
	hps_hps_io_hps_io_emac1_inst_RXD3,
	hps_hps_io_hps_io_sdio_inst_CMD,
	hps_hps_io_hps_io_sdio_inst_D0,
	hps_hps_io_hps_io_sdio_inst_D1,
	hps_hps_io_hps_io_sdio_inst_CLK,
	hps_hps_io_hps_io_sdio_inst_D2,
	hps_hps_io_hps_io_sdio_inst_D3,
	hps_hps_io_hps_io_uart0_inst_RX,
	hps_hps_io_hps_io_uart0_inst_TX,
	leds_out_export,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	reset_reset_n,
	state_in_export,
	switches_in_export)/* synthesis synthesis_greybox=0 */;
output 	[31:0] base_addr_ddr_out_export;
input 	clk_clk;
output 	[31:0] control_out_export;
input 	[26:0] hps_f2h_sdram0_data_address;
input 	[7:0] hps_f2h_sdram0_data_burstcount;
output 	hps_f2h_sdram0_data_waitrequest;
output 	[255:0] hps_f2h_sdram0_data_readdata;
output 	hps_f2h_sdram0_data_readdatavalid;
input 	hps_f2h_sdram0_data_read;
input 	[255:0] hps_f2h_sdram0_data_writedata;
input 	[31:0] hps_f2h_sdram0_data_byteenable;
input 	hps_f2h_sdram0_data_write;
input 	[27:0] hps_f2h_stm_hw_events_stm_hwevents;
output 	hps_h2f_cold_reset_reset_n;
output 	hps_h2f_warm_reset_handshake_h2f_pending_rst_req_n;
input 	hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n;
output 	hps_hps_io_hps_io_emac1_inst_TX_CLK;
output 	hps_hps_io_hps_io_emac1_inst_TXD0;
output 	hps_hps_io_hps_io_emac1_inst_TXD1;
output 	hps_hps_io_hps_io_emac1_inst_TXD2;
output 	hps_hps_io_hps_io_emac1_inst_TXD3;
input 	hps_hps_io_hps_io_emac1_inst_RXD0;
inout 	hps_hps_io_hps_io_emac1_inst_MDIO;
output 	hps_hps_io_hps_io_emac1_inst_MDC;
input 	hps_hps_io_hps_io_emac1_inst_RX_CTL;
output 	hps_hps_io_hps_io_emac1_inst_TX_CTL;
input 	hps_hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_hps_io_hps_io_emac1_inst_RXD1;
input 	hps_hps_io_hps_io_emac1_inst_RXD2;
input 	hps_hps_io_hps_io_emac1_inst_RXD3;
inout 	hps_hps_io_hps_io_sdio_inst_CMD;
inout 	hps_hps_io_hps_io_sdio_inst_D0;
inout 	hps_hps_io_hps_io_sdio_inst_D1;
output 	hps_hps_io_hps_io_sdio_inst_CLK;
inout 	hps_hps_io_hps_io_sdio_inst_D2;
inout 	hps_hps_io_hps_io_sdio_inst_D3;
input 	hps_hps_io_hps_io_uart0_inst_RX;
output 	hps_hps_io_hps_io_uart0_inst_TX;
output 	[9:0] leds_out_export;
output 	[14:0] memory_mem_a;
output 	[2:0] memory_mem_ba;
output 	memory_mem_ck;
output 	memory_mem_ck_n;
output 	memory_mem_cke;
output 	memory_mem_cs_n;
output 	memory_mem_ras_n;
output 	memory_mem_cas_n;
output 	memory_mem_we_n;
output 	memory_mem_reset_n;
inout 	[31:0] memory_mem_dq;
inout 	[3:0] memory_mem_dqs;
inout 	[3:0] memory_mem_dqs_n;
output 	memory_mem_odt;
output 	[3:0] memory_mem_dm;
input 	memory_oct_rzqin;
input 	reset_reset_n;
input 	[31:0] state_in_export;
input 	[9:0] switches_in_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps|fpga_interfaces|h2f_cold_rst_n[0] ;
wire \hps|fpga_interfaces|h2f_pending_rst_req_n[0] ;
wire \hps|fpga_interfaces|h2f_rst_n[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARVALID[0] ;
wire \hps|fpga_interfaces|h2f_lw_AWVALID[0] ;
wire \hps|fpga_interfaces|h2f_lw_BREADY[0] ;
wire \hps|fpga_interfaces|h2f_lw_RREADY[0] ;
wire \hps|fpga_interfaces|h2f_lw_WLAST[0] ;
wire \hps|fpga_interfaces|h2f_lw_WVALID[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[1] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[2] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[3] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[4] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[5] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[6] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[7] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[8] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[9] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[10] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[11] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[12] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[13] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[14] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[15] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[16] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[17] ;
wire \hps|fpga_interfaces|h2f_lw_ARADDR[18] ;
wire \hps|fpga_interfaces|h2f_lw_ARBURST[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARBURST[1] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[1] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[2] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[3] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[4] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[5] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[6] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[7] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[8] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[9] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[10] ;
wire \hps|fpga_interfaces|h2f_lw_ARID[11] ;
wire \hps|fpga_interfaces|h2f_lw_ARLEN[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARLEN[1] ;
wire \hps|fpga_interfaces|h2f_lw_ARLEN[2] ;
wire \hps|fpga_interfaces|h2f_lw_ARLEN[3] ;
wire \hps|fpga_interfaces|h2f_lw_ARSIZE[0] ;
wire \hps|fpga_interfaces|h2f_lw_ARSIZE[1] ;
wire \hps|fpga_interfaces|h2f_lw_ARSIZE[2] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[0] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[1] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[2] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[3] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[4] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[5] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[6] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[7] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[8] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[9] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[10] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[11] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[12] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[13] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[14] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[15] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[16] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[17] ;
wire \hps|fpga_interfaces|h2f_lw_AWADDR[18] ;
wire \hps|fpga_interfaces|h2f_lw_AWBURST[0] ;
wire \hps|fpga_interfaces|h2f_lw_AWBURST[1] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[0] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[1] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[2] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[3] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[4] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[5] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[6] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[7] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[8] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[9] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[10] ;
wire \hps|fpga_interfaces|h2f_lw_AWID[11] ;
wire \hps|fpga_interfaces|h2f_lw_AWLEN[0] ;
wire \hps|fpga_interfaces|h2f_lw_AWLEN[1] ;
wire \hps|fpga_interfaces|h2f_lw_AWLEN[2] ;
wire \hps|fpga_interfaces|h2f_lw_AWLEN[3] ;
wire \hps|fpga_interfaces|h2f_lw_AWSIZE[0] ;
wire \hps|fpga_interfaces|h2f_lw_AWSIZE[1] ;
wire \hps|fpga_interfaces|h2f_lw_AWSIZE[2] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[0] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[1] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[2] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[3] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[4] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[5] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[6] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[7] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[8] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[9] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[10] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[11] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[12] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[13] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[14] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[15] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[16] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[17] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[18] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[19] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[20] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[21] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[22] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[23] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[24] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[25] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[26] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[27] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[28] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[29] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[30] ;
wire \hps|fpga_interfaces|h2f_lw_WDATA[31] ;
wire \hps|fpga_interfaces|h2f_lw_WSTRB[0] ;
wire \hps|fpga_interfaces|h2f_lw_WSTRB[1] ;
wire \hps|fpga_interfaces|h2f_lw_WSTRB[2] ;
wire \hps|fpga_interfaces|h2f_lw_WSTRB[3] ;
wire \hps|fpga_interfaces|intermediate[1] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATAVALID[0] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[0] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[1] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[2] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[3] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[4] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[5] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[6] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[7] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[8] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[9] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[10] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[11] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[12] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[13] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[14] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[15] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[16] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[17] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[18] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[19] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[20] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[21] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[22] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[23] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[24] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[25] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[26] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[27] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[28] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[29] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[30] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[31] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[32] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[33] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[34] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[35] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[36] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[37] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[38] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[39] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[40] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[41] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[42] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[43] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[44] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[45] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[46] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[47] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[48] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[49] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[50] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[51] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[52] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[53] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[54] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[55] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[56] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[57] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[58] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[59] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[60] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[61] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[62] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[63] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[64] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[65] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[66] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[67] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[68] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[69] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[70] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[71] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[72] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[73] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[74] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[75] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[76] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[77] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[78] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[79] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[80] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[81] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[82] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[83] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[84] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[85] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[86] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[87] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[88] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[89] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[90] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[91] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[92] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[93] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[94] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[95] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[96] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[97] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[98] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[99] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[100] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[101] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[102] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[103] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[104] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[105] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[106] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[107] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[108] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[109] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[110] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[111] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[112] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[113] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[114] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[115] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[116] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[117] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[118] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[119] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[120] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[121] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[122] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[123] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[124] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[125] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[126] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[127] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[128] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[129] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[130] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[131] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[132] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[133] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[134] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[135] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[136] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[137] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[138] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[139] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[140] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[141] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[142] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[143] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[144] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[145] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[146] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[147] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[148] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[149] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[150] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[151] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[152] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[153] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[154] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[155] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[156] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[157] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[158] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[159] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[160] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[161] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[162] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[163] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[164] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[165] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[166] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[167] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[168] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[169] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[170] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[171] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[172] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[173] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[174] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[175] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[176] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[177] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[178] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[179] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[180] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[181] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[182] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[183] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[184] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[185] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[186] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[187] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[188] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[189] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[190] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[191] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[192] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[193] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[194] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[195] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[196] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[197] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[198] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[199] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[200] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[201] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[202] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[203] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[204] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[205] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[206] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[207] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[208] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[209] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[210] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[211] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[212] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[213] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[214] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[215] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[216] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[217] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[218] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[219] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[220] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[221] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[222] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[223] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[224] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[225] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[226] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[227] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[228] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[229] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[230] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[231] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[232] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[233] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[234] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[235] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[236] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[237] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[238] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[239] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[240] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[241] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[242] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[243] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[244] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[245] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[246] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[247] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[248] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[249] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[250] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[251] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[252] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[253] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[254] ;
wire \hps|fpga_interfaces|f2h_sdram0_READDATA[255] ;
wire \base_address_ddr|data_out[0]~q ;
wire \base_address_ddr|data_out[1]~q ;
wire \base_address_ddr|data_out[2]~q ;
wire \base_address_ddr|data_out[3]~q ;
wire \base_address_ddr|data_out[4]~q ;
wire \base_address_ddr|data_out[5]~q ;
wire \base_address_ddr|data_out[6]~q ;
wire \base_address_ddr|data_out[7]~q ;
wire \base_address_ddr|data_out[8]~q ;
wire \base_address_ddr|data_out[9]~q ;
wire \base_address_ddr|data_out[10]~q ;
wire \base_address_ddr|data_out[11]~q ;
wire \base_address_ddr|data_out[12]~q ;
wire \base_address_ddr|data_out[13]~q ;
wire \base_address_ddr|data_out[14]~q ;
wire \base_address_ddr|data_out[15]~q ;
wire \base_address_ddr|data_out[16]~q ;
wire \base_address_ddr|data_out[17]~q ;
wire \base_address_ddr|data_out[18]~q ;
wire \base_address_ddr|data_out[19]~q ;
wire \base_address_ddr|data_out[20]~q ;
wire \base_address_ddr|data_out[21]~q ;
wire \base_address_ddr|data_out[22]~q ;
wire \base_address_ddr|data_out[23]~q ;
wire \base_address_ddr|data_out[24]~q ;
wire \base_address_ddr|data_out[25]~q ;
wire \base_address_ddr|data_out[26]~q ;
wire \base_address_ddr|data_out[27]~q ;
wire \base_address_ddr|data_out[28]~q ;
wire \base_address_ddr|data_out[29]~q ;
wire \base_address_ddr|data_out[30]~q ;
wire \base_address_ddr|data_out[31]~q ;
wire \control|data_out[0]~q ;
wire \control|data_out[1]~q ;
wire \control|data_out[2]~q ;
wire \control|data_out[3]~q ;
wire \control|data_out[4]~q ;
wire \control|data_out[5]~q ;
wire \control|data_out[6]~q ;
wire \control|data_out[7]~q ;
wire \control|data_out[8]~q ;
wire \control|data_out[9]~q ;
wire \control|data_out[10]~q ;
wire \control|data_out[11]~q ;
wire \control|data_out[12]~q ;
wire \control|data_out[13]~q ;
wire \control|data_out[14]~q ;
wire \control|data_out[15]~q ;
wire \control|data_out[16]~q ;
wire \control|data_out[17]~q ;
wire \control|data_out[18]~q ;
wire \control|data_out[19]~q ;
wire \control|data_out[20]~q ;
wire \control|data_out[21]~q ;
wire \control|data_out[22]~q ;
wire \control|data_out[23]~q ;
wire \control|data_out[24]~q ;
wire \control|data_out[25]~q ;
wire \control|data_out[26]~q ;
wire \control|data_out[27]~q ;
wire \control|data_out[28]~q ;
wire \control|data_out[29]~q ;
wire \control|data_out[30]~q ;
wire \control|data_out[31]~q ;
wire \leds|data_out[0]~q ;
wire \leds|data_out[1]~q ;
wire \leds|data_out[2]~q ;
wire \leds|data_out[3]~q ;
wire \leds|data_out[4]~q ;
wire \leds|data_out[5]~q ;
wire \leds|data_out[6]~q ;
wire \leds|data_out[7]~q ;
wire \leds|data_out[8]~q ;
wire \leds|data_out[9]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|control_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|control_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|leds_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|leds_s1_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|hps_h2f_lw_axi_master_rd_limiter|cmd_sink_ready~0_combout ;
wire \mm_interconnect_0|hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~2_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~3_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~4_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~5_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~6_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~7_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~8_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~9_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~10_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~11_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~5_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[1]~11_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~17_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~23_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[4]~29_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~35_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~41_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~48_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~54_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~58_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~11_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~14_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~17_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~20_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~23_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~26_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~29_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~32_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~35_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~38_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~41_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~44_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~47_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~50_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~53_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~56_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~59_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~62_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~65_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~68_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~71_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_payload~74_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[92]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[93]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[94]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[95]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[96]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[97]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[98]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[99]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[100]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[101]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[102]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[103]~combout ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \rst_controller|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|base_address_ddr_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \rst_controller_001|rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \mm_interconnect_0|control_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ;
wire \mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ;
wire \mm_interconnect_0|leds_s1_agent|m0_write~combout ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ;
wire \mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ;
wire \rst_controller_002|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \control|readdata[0]~combout ;
wire \base_address_ddr|readdata[0]~combout ;
wire \leds|readdata[0]~combout ;
wire \state|readdata[0]~q ;
wire \switches|readdata[0]~q ;
wire \control|readdata[1]~combout ;
wire \base_address_ddr|readdata[1]~combout ;
wire \leds|readdata[1]~combout ;
wire \state|readdata[1]~q ;
wire \switches|readdata[1]~q ;
wire \control|readdata[2]~combout ;
wire \base_address_ddr|readdata[2]~combout ;
wire \leds|readdata[2]~combout ;
wire \state|readdata[2]~q ;
wire \switches|readdata[2]~q ;
wire \control|readdata[3]~combout ;
wire \base_address_ddr|readdata[3]~combout ;
wire \leds|readdata[3]~combout ;
wire \state|readdata[3]~q ;
wire \switches|readdata[3]~q ;
wire \control|readdata[4]~combout ;
wire \base_address_ddr|readdata[4]~combout ;
wire \leds|readdata[4]~combout ;
wire \state|readdata[4]~q ;
wire \switches|readdata[4]~q ;
wire \control|readdata[5]~combout ;
wire \base_address_ddr|readdata[5]~combout ;
wire \leds|readdata[5]~combout ;
wire \state|readdata[5]~q ;
wire \switches|readdata[5]~q ;
wire \control|readdata[6]~combout ;
wire \base_address_ddr|readdata[6]~combout ;
wire \leds|readdata[6]~combout ;
wire \state|readdata[6]~q ;
wire \switches|readdata[6]~q ;
wire \control|readdata[7]~combout ;
wire \base_address_ddr|readdata[7]~combout ;
wire \leds|readdata[7]~combout ;
wire \state|readdata[7]~q ;
wire \switches|readdata[7]~q ;
wire \control|readdata[8]~combout ;
wire \base_address_ddr|readdata[8]~combout ;
wire \leds|readdata[8]~combout ;
wire \state|readdata[8]~q ;
wire \switches|readdata[8]~q ;
wire \state|readdata[9]~q ;
wire \control|readdata[9]~combout ;
wire \base_address_ddr|readdata[9]~combout ;
wire \leds|readdata[9]~combout ;
wire \switches|readdata[9]~q ;
wire \control|readdata[10]~combout ;
wire \base_address_ddr|readdata[10]~combout ;
wire \state|readdata[10]~q ;
wire \control|readdata[11]~combout ;
wire \base_address_ddr|readdata[11]~combout ;
wire \state|readdata[11]~q ;
wire \base_address_ddr|readdata[12]~combout ;
wire \control|readdata[12]~combout ;
wire \state|readdata[12]~q ;
wire \base_address_ddr|readdata[13]~combout ;
wire \control|readdata[13]~combout ;
wire \state|readdata[13]~q ;
wire \base_address_ddr|readdata[14]~combout ;
wire \control|readdata[14]~combout ;
wire \state|readdata[14]~q ;
wire \base_address_ddr|readdata[15]~combout ;
wire \control|readdata[15]~combout ;
wire \state|readdata[15]~q ;
wire \base_address_ddr|readdata[16]~combout ;
wire \control|readdata[16]~combout ;
wire \state|readdata[16]~q ;
wire \base_address_ddr|readdata[17]~combout ;
wire \control|readdata[17]~combout ;
wire \state|readdata[17]~q ;
wire \base_address_ddr|readdata[18]~combout ;
wire \control|readdata[18]~combout ;
wire \state|readdata[18]~q ;
wire \control|readdata[19]~combout ;
wire \base_address_ddr|readdata[19]~combout ;
wire \state|readdata[19]~q ;
wire \control|readdata[20]~combout ;
wire \base_address_ddr|readdata[20]~combout ;
wire \state|readdata[20]~q ;
wire \control|readdata[21]~combout ;
wire \base_address_ddr|readdata[21]~combout ;
wire \state|readdata[21]~q ;
wire \base_address_ddr|readdata[22]~combout ;
wire \control|readdata[22]~combout ;
wire \state|readdata[22]~q ;
wire \base_address_ddr|readdata[23]~combout ;
wire \control|readdata[23]~combout ;
wire \state|readdata[23]~q ;
wire \control|readdata[24]~combout ;
wire \base_address_ddr|readdata[24]~combout ;
wire \state|readdata[24]~q ;
wire \base_address_ddr|readdata[25]~combout ;
wire \control|readdata[25]~combout ;
wire \state|readdata[25]~q ;
wire \base_address_ddr|readdata[26]~combout ;
wire \control|readdata[26]~combout ;
wire \state|readdata[26]~q ;
wire \control|readdata[27]~combout ;
wire \base_address_ddr|readdata[27]~combout ;
wire \state|readdata[27]~q ;
wire \control|readdata[28]~combout ;
wire \base_address_ddr|readdata[28]~combout ;
wire \state|readdata[28]~q ;
wire \base_address_ddr|readdata[29]~combout ;
wire \control|readdata[29]~combout ;
wire \state|readdata[29]~q ;
wire \control|readdata[30]~combout ;
wire \base_address_ddr|readdata[30]~combout ;
wire \state|readdata[30]~q ;
wire \base_address_ddr|readdata[31]~combout ;
wire \control|readdata[31]~combout ;
wire \state|readdata[31]~q ;
wire \mm_interconnect_0|state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \mm_interconnect_0|switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ;
wire \mm_interconnect_0|switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;
wire \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;
wire \hps|hps_io|border|intermediate[0] ;
wire \hps|hps_io|border|intermediate[1] ;
wire \hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;
wire \hps|hps_io|border|emac1_inst~emac_phy_txd ;
wire \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;
wire \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;
wire \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;
wire \hps|hps_io|border|sdio_inst~sdmmc_cclk ;
wire \hps|hps_io|border|intermediate[2] ;
wire \hps|hps_io|border|intermediate[3] ;
wire \hps|hps_io|border|intermediate[4] ;
wire \hps|hps_io|border|intermediate[6] ;
wire \hps|hps_io|border|intermediate[8] ;
wire \hps|hps_io|border|intermediate[10] ;
wire \hps|hps_io|border|intermediate[5] ;
wire \hps|hps_io|border|intermediate[7] ;
wire \hps|hps_io|border|intermediate[9] ;
wire \hps|hps_io|border|intermediate[11] ;
wire \hps|hps_io|border|uart0_inst~uart_txd ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ;
wire \hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ;
wire \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ;
wire \hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ;
wire \hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ;
wire \hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ;
wire \hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ;
wire \hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ;
wire \hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[0]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[1]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[2]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[3]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[4]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[5]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[6]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[7]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[8]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[9]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[10]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[11]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[12]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[13]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[14]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[15]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[16]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[17]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[18]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[19]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[20]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[21]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[22]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[23]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[24]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[25]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[26]~input_o ;
wire \hps_f2h_stm_hw_events_stm_hwevents[27]~input_o ;
wire \clk_clk~input_o ;
wire \hps_hps_io_hps_io_emac1_inst_RXD0~input_o ;
wire \hps_hps_io_hps_io_emac1_inst_RXD1~input_o ;
wire \hps_hps_io_hps_io_emac1_inst_RXD2~input_o ;
wire \hps_hps_io_hps_io_emac1_inst_RXD3~input_o ;
wire \hps_hps_io_hps_io_emac1_inst_RX_CLK~input_o ;
wire \hps_hps_io_hps_io_emac1_inst_RX_CTL~input_o ;
wire \hps_hps_io_hps_io_uart0_inst_RX~input_o ;
wire \memory_oct_rzqin~input_o ;
wire \hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n~input_o ;
wire \hps_f2h_sdram0_data_read~input_o ;
wire \hps_f2h_sdram0_data_write~input_o ;
wire \hps_f2h_sdram0_data_address[0]~input_o ;
wire \hps_f2h_sdram0_data_address[1]~input_o ;
wire \hps_f2h_sdram0_data_address[2]~input_o ;
wire \hps_f2h_sdram0_data_address[3]~input_o ;
wire \hps_f2h_sdram0_data_address[4]~input_o ;
wire \hps_f2h_sdram0_data_address[5]~input_o ;
wire \hps_f2h_sdram0_data_address[6]~input_o ;
wire \hps_f2h_sdram0_data_address[7]~input_o ;
wire \hps_f2h_sdram0_data_address[8]~input_o ;
wire \hps_f2h_sdram0_data_address[9]~input_o ;
wire \hps_f2h_sdram0_data_address[10]~input_o ;
wire \hps_f2h_sdram0_data_address[11]~input_o ;
wire \hps_f2h_sdram0_data_address[12]~input_o ;
wire \hps_f2h_sdram0_data_address[13]~input_o ;
wire \hps_f2h_sdram0_data_address[14]~input_o ;
wire \hps_f2h_sdram0_data_address[15]~input_o ;
wire \hps_f2h_sdram0_data_address[16]~input_o ;
wire \hps_f2h_sdram0_data_address[17]~input_o ;
wire \hps_f2h_sdram0_data_address[18]~input_o ;
wire \hps_f2h_sdram0_data_address[19]~input_o ;
wire \hps_f2h_sdram0_data_address[20]~input_o ;
wire \hps_f2h_sdram0_data_address[21]~input_o ;
wire \hps_f2h_sdram0_data_address[22]~input_o ;
wire \hps_f2h_sdram0_data_address[23]~input_o ;
wire \hps_f2h_sdram0_data_address[24]~input_o ;
wire \hps_f2h_sdram0_data_address[25]~input_o ;
wire \hps_f2h_sdram0_data_address[26]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[0]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[1]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[2]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[3]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[4]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[5]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[6]~input_o ;
wire \hps_f2h_sdram0_data_burstcount[7]~input_o ;
wire \hps_f2h_sdram0_data_writedata[0]~input_o ;
wire \hps_f2h_sdram0_data_writedata[1]~input_o ;
wire \hps_f2h_sdram0_data_writedata[2]~input_o ;
wire \hps_f2h_sdram0_data_writedata[3]~input_o ;
wire \hps_f2h_sdram0_data_writedata[4]~input_o ;
wire \hps_f2h_sdram0_data_writedata[5]~input_o ;
wire \hps_f2h_sdram0_data_writedata[6]~input_o ;
wire \hps_f2h_sdram0_data_writedata[7]~input_o ;
wire \hps_f2h_sdram0_data_writedata[8]~input_o ;
wire \hps_f2h_sdram0_data_writedata[9]~input_o ;
wire \hps_f2h_sdram0_data_writedata[10]~input_o ;
wire \hps_f2h_sdram0_data_writedata[11]~input_o ;
wire \hps_f2h_sdram0_data_writedata[12]~input_o ;
wire \hps_f2h_sdram0_data_writedata[13]~input_o ;
wire \hps_f2h_sdram0_data_writedata[14]~input_o ;
wire \hps_f2h_sdram0_data_writedata[15]~input_o ;
wire \hps_f2h_sdram0_data_writedata[16]~input_o ;
wire \hps_f2h_sdram0_data_writedata[17]~input_o ;
wire \hps_f2h_sdram0_data_writedata[18]~input_o ;
wire \hps_f2h_sdram0_data_writedata[19]~input_o ;
wire \hps_f2h_sdram0_data_writedata[20]~input_o ;
wire \hps_f2h_sdram0_data_writedata[21]~input_o ;
wire \hps_f2h_sdram0_data_writedata[22]~input_o ;
wire \hps_f2h_sdram0_data_writedata[23]~input_o ;
wire \hps_f2h_sdram0_data_writedata[24]~input_o ;
wire \hps_f2h_sdram0_data_writedata[25]~input_o ;
wire \hps_f2h_sdram0_data_writedata[26]~input_o ;
wire \hps_f2h_sdram0_data_writedata[27]~input_o ;
wire \hps_f2h_sdram0_data_writedata[28]~input_o ;
wire \hps_f2h_sdram0_data_writedata[29]~input_o ;
wire \hps_f2h_sdram0_data_writedata[30]~input_o ;
wire \hps_f2h_sdram0_data_writedata[31]~input_o ;
wire \hps_f2h_sdram0_data_writedata[32]~input_o ;
wire \hps_f2h_sdram0_data_writedata[33]~input_o ;
wire \hps_f2h_sdram0_data_writedata[34]~input_o ;
wire \hps_f2h_sdram0_data_writedata[35]~input_o ;
wire \hps_f2h_sdram0_data_writedata[36]~input_o ;
wire \hps_f2h_sdram0_data_writedata[37]~input_o ;
wire \hps_f2h_sdram0_data_writedata[38]~input_o ;
wire \hps_f2h_sdram0_data_writedata[39]~input_o ;
wire \hps_f2h_sdram0_data_writedata[40]~input_o ;
wire \hps_f2h_sdram0_data_writedata[41]~input_o ;
wire \hps_f2h_sdram0_data_writedata[42]~input_o ;
wire \hps_f2h_sdram0_data_writedata[43]~input_o ;
wire \hps_f2h_sdram0_data_writedata[44]~input_o ;
wire \hps_f2h_sdram0_data_writedata[45]~input_o ;
wire \hps_f2h_sdram0_data_writedata[46]~input_o ;
wire \hps_f2h_sdram0_data_writedata[47]~input_o ;
wire \hps_f2h_sdram0_data_writedata[48]~input_o ;
wire \hps_f2h_sdram0_data_writedata[49]~input_o ;
wire \hps_f2h_sdram0_data_writedata[50]~input_o ;
wire \hps_f2h_sdram0_data_writedata[51]~input_o ;
wire \hps_f2h_sdram0_data_writedata[52]~input_o ;
wire \hps_f2h_sdram0_data_writedata[53]~input_o ;
wire \hps_f2h_sdram0_data_writedata[54]~input_o ;
wire \hps_f2h_sdram0_data_writedata[55]~input_o ;
wire \hps_f2h_sdram0_data_writedata[56]~input_o ;
wire \hps_f2h_sdram0_data_writedata[57]~input_o ;
wire \hps_f2h_sdram0_data_writedata[58]~input_o ;
wire \hps_f2h_sdram0_data_writedata[59]~input_o ;
wire \hps_f2h_sdram0_data_writedata[60]~input_o ;
wire \hps_f2h_sdram0_data_writedata[61]~input_o ;
wire \hps_f2h_sdram0_data_writedata[62]~input_o ;
wire \hps_f2h_sdram0_data_writedata[63]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[0]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[1]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[2]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[3]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[4]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[5]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[6]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[7]~input_o ;
wire \hps_f2h_sdram0_data_writedata[64]~input_o ;
wire \hps_f2h_sdram0_data_writedata[65]~input_o ;
wire \hps_f2h_sdram0_data_writedata[66]~input_o ;
wire \hps_f2h_sdram0_data_writedata[67]~input_o ;
wire \hps_f2h_sdram0_data_writedata[68]~input_o ;
wire \hps_f2h_sdram0_data_writedata[69]~input_o ;
wire \hps_f2h_sdram0_data_writedata[70]~input_o ;
wire \hps_f2h_sdram0_data_writedata[71]~input_o ;
wire \hps_f2h_sdram0_data_writedata[72]~input_o ;
wire \hps_f2h_sdram0_data_writedata[73]~input_o ;
wire \hps_f2h_sdram0_data_writedata[74]~input_o ;
wire \hps_f2h_sdram0_data_writedata[75]~input_o ;
wire \hps_f2h_sdram0_data_writedata[76]~input_o ;
wire \hps_f2h_sdram0_data_writedata[77]~input_o ;
wire \hps_f2h_sdram0_data_writedata[78]~input_o ;
wire \hps_f2h_sdram0_data_writedata[79]~input_o ;
wire \hps_f2h_sdram0_data_writedata[80]~input_o ;
wire \hps_f2h_sdram0_data_writedata[81]~input_o ;
wire \hps_f2h_sdram0_data_writedata[82]~input_o ;
wire \hps_f2h_sdram0_data_writedata[83]~input_o ;
wire \hps_f2h_sdram0_data_writedata[84]~input_o ;
wire \hps_f2h_sdram0_data_writedata[85]~input_o ;
wire \hps_f2h_sdram0_data_writedata[86]~input_o ;
wire \hps_f2h_sdram0_data_writedata[87]~input_o ;
wire \hps_f2h_sdram0_data_writedata[88]~input_o ;
wire \hps_f2h_sdram0_data_writedata[89]~input_o ;
wire \hps_f2h_sdram0_data_writedata[90]~input_o ;
wire \hps_f2h_sdram0_data_writedata[91]~input_o ;
wire \hps_f2h_sdram0_data_writedata[92]~input_o ;
wire \hps_f2h_sdram0_data_writedata[93]~input_o ;
wire \hps_f2h_sdram0_data_writedata[94]~input_o ;
wire \hps_f2h_sdram0_data_writedata[95]~input_o ;
wire \hps_f2h_sdram0_data_writedata[96]~input_o ;
wire \hps_f2h_sdram0_data_writedata[97]~input_o ;
wire \hps_f2h_sdram0_data_writedata[98]~input_o ;
wire \hps_f2h_sdram0_data_writedata[99]~input_o ;
wire \hps_f2h_sdram0_data_writedata[100]~input_o ;
wire \hps_f2h_sdram0_data_writedata[101]~input_o ;
wire \hps_f2h_sdram0_data_writedata[102]~input_o ;
wire \hps_f2h_sdram0_data_writedata[103]~input_o ;
wire \hps_f2h_sdram0_data_writedata[104]~input_o ;
wire \hps_f2h_sdram0_data_writedata[105]~input_o ;
wire \hps_f2h_sdram0_data_writedata[106]~input_o ;
wire \hps_f2h_sdram0_data_writedata[107]~input_o ;
wire \hps_f2h_sdram0_data_writedata[108]~input_o ;
wire \hps_f2h_sdram0_data_writedata[109]~input_o ;
wire \hps_f2h_sdram0_data_writedata[110]~input_o ;
wire \hps_f2h_sdram0_data_writedata[111]~input_o ;
wire \hps_f2h_sdram0_data_writedata[112]~input_o ;
wire \hps_f2h_sdram0_data_writedata[113]~input_o ;
wire \hps_f2h_sdram0_data_writedata[114]~input_o ;
wire \hps_f2h_sdram0_data_writedata[115]~input_o ;
wire \hps_f2h_sdram0_data_writedata[116]~input_o ;
wire \hps_f2h_sdram0_data_writedata[117]~input_o ;
wire \hps_f2h_sdram0_data_writedata[118]~input_o ;
wire \hps_f2h_sdram0_data_writedata[119]~input_o ;
wire \hps_f2h_sdram0_data_writedata[120]~input_o ;
wire \hps_f2h_sdram0_data_writedata[121]~input_o ;
wire \hps_f2h_sdram0_data_writedata[122]~input_o ;
wire \hps_f2h_sdram0_data_writedata[123]~input_o ;
wire \hps_f2h_sdram0_data_writedata[124]~input_o ;
wire \hps_f2h_sdram0_data_writedata[125]~input_o ;
wire \hps_f2h_sdram0_data_writedata[126]~input_o ;
wire \hps_f2h_sdram0_data_writedata[127]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[8]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[9]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[10]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[11]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[12]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[13]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[14]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[15]~input_o ;
wire \hps_f2h_sdram0_data_writedata[128]~input_o ;
wire \hps_f2h_sdram0_data_writedata[129]~input_o ;
wire \hps_f2h_sdram0_data_writedata[130]~input_o ;
wire \hps_f2h_sdram0_data_writedata[131]~input_o ;
wire \hps_f2h_sdram0_data_writedata[132]~input_o ;
wire \hps_f2h_sdram0_data_writedata[133]~input_o ;
wire \hps_f2h_sdram0_data_writedata[134]~input_o ;
wire \hps_f2h_sdram0_data_writedata[135]~input_o ;
wire \hps_f2h_sdram0_data_writedata[136]~input_o ;
wire \hps_f2h_sdram0_data_writedata[137]~input_o ;
wire \hps_f2h_sdram0_data_writedata[138]~input_o ;
wire \hps_f2h_sdram0_data_writedata[139]~input_o ;
wire \hps_f2h_sdram0_data_writedata[140]~input_o ;
wire \hps_f2h_sdram0_data_writedata[141]~input_o ;
wire \hps_f2h_sdram0_data_writedata[142]~input_o ;
wire \hps_f2h_sdram0_data_writedata[143]~input_o ;
wire \hps_f2h_sdram0_data_writedata[144]~input_o ;
wire \hps_f2h_sdram0_data_writedata[145]~input_o ;
wire \hps_f2h_sdram0_data_writedata[146]~input_o ;
wire \hps_f2h_sdram0_data_writedata[147]~input_o ;
wire \hps_f2h_sdram0_data_writedata[148]~input_o ;
wire \hps_f2h_sdram0_data_writedata[149]~input_o ;
wire \hps_f2h_sdram0_data_writedata[150]~input_o ;
wire \hps_f2h_sdram0_data_writedata[151]~input_o ;
wire \hps_f2h_sdram0_data_writedata[152]~input_o ;
wire \hps_f2h_sdram0_data_writedata[153]~input_o ;
wire \hps_f2h_sdram0_data_writedata[154]~input_o ;
wire \hps_f2h_sdram0_data_writedata[155]~input_o ;
wire \hps_f2h_sdram0_data_writedata[156]~input_o ;
wire \hps_f2h_sdram0_data_writedata[157]~input_o ;
wire \hps_f2h_sdram0_data_writedata[158]~input_o ;
wire \hps_f2h_sdram0_data_writedata[159]~input_o ;
wire \hps_f2h_sdram0_data_writedata[160]~input_o ;
wire \hps_f2h_sdram0_data_writedata[161]~input_o ;
wire \hps_f2h_sdram0_data_writedata[162]~input_o ;
wire \hps_f2h_sdram0_data_writedata[163]~input_o ;
wire \hps_f2h_sdram0_data_writedata[164]~input_o ;
wire \hps_f2h_sdram0_data_writedata[165]~input_o ;
wire \hps_f2h_sdram0_data_writedata[166]~input_o ;
wire \hps_f2h_sdram0_data_writedata[167]~input_o ;
wire \hps_f2h_sdram0_data_writedata[168]~input_o ;
wire \hps_f2h_sdram0_data_writedata[169]~input_o ;
wire \hps_f2h_sdram0_data_writedata[170]~input_o ;
wire \hps_f2h_sdram0_data_writedata[171]~input_o ;
wire \hps_f2h_sdram0_data_writedata[172]~input_o ;
wire \hps_f2h_sdram0_data_writedata[173]~input_o ;
wire \hps_f2h_sdram0_data_writedata[174]~input_o ;
wire \hps_f2h_sdram0_data_writedata[175]~input_o ;
wire \hps_f2h_sdram0_data_writedata[176]~input_o ;
wire \hps_f2h_sdram0_data_writedata[177]~input_o ;
wire \hps_f2h_sdram0_data_writedata[178]~input_o ;
wire \hps_f2h_sdram0_data_writedata[179]~input_o ;
wire \hps_f2h_sdram0_data_writedata[180]~input_o ;
wire \hps_f2h_sdram0_data_writedata[181]~input_o ;
wire \hps_f2h_sdram0_data_writedata[182]~input_o ;
wire \hps_f2h_sdram0_data_writedata[183]~input_o ;
wire \hps_f2h_sdram0_data_writedata[184]~input_o ;
wire \hps_f2h_sdram0_data_writedata[185]~input_o ;
wire \hps_f2h_sdram0_data_writedata[186]~input_o ;
wire \hps_f2h_sdram0_data_writedata[187]~input_o ;
wire \hps_f2h_sdram0_data_writedata[188]~input_o ;
wire \hps_f2h_sdram0_data_writedata[189]~input_o ;
wire \hps_f2h_sdram0_data_writedata[190]~input_o ;
wire \hps_f2h_sdram0_data_writedata[191]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[16]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[17]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[18]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[19]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[20]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[21]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[22]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[23]~input_o ;
wire \hps_f2h_sdram0_data_writedata[192]~input_o ;
wire \hps_f2h_sdram0_data_writedata[193]~input_o ;
wire \hps_f2h_sdram0_data_writedata[194]~input_o ;
wire \hps_f2h_sdram0_data_writedata[195]~input_o ;
wire \hps_f2h_sdram0_data_writedata[196]~input_o ;
wire \hps_f2h_sdram0_data_writedata[197]~input_o ;
wire \hps_f2h_sdram0_data_writedata[198]~input_o ;
wire \hps_f2h_sdram0_data_writedata[199]~input_o ;
wire \hps_f2h_sdram0_data_writedata[200]~input_o ;
wire \hps_f2h_sdram0_data_writedata[201]~input_o ;
wire \hps_f2h_sdram0_data_writedata[202]~input_o ;
wire \hps_f2h_sdram0_data_writedata[203]~input_o ;
wire \hps_f2h_sdram0_data_writedata[204]~input_o ;
wire \hps_f2h_sdram0_data_writedata[205]~input_o ;
wire \hps_f2h_sdram0_data_writedata[206]~input_o ;
wire \hps_f2h_sdram0_data_writedata[207]~input_o ;
wire \hps_f2h_sdram0_data_writedata[208]~input_o ;
wire \hps_f2h_sdram0_data_writedata[209]~input_o ;
wire \hps_f2h_sdram0_data_writedata[210]~input_o ;
wire \hps_f2h_sdram0_data_writedata[211]~input_o ;
wire \hps_f2h_sdram0_data_writedata[212]~input_o ;
wire \hps_f2h_sdram0_data_writedata[213]~input_o ;
wire \hps_f2h_sdram0_data_writedata[214]~input_o ;
wire \hps_f2h_sdram0_data_writedata[215]~input_o ;
wire \hps_f2h_sdram0_data_writedata[216]~input_o ;
wire \hps_f2h_sdram0_data_writedata[217]~input_o ;
wire \hps_f2h_sdram0_data_writedata[218]~input_o ;
wire \hps_f2h_sdram0_data_writedata[219]~input_o ;
wire \hps_f2h_sdram0_data_writedata[220]~input_o ;
wire \hps_f2h_sdram0_data_writedata[221]~input_o ;
wire \hps_f2h_sdram0_data_writedata[222]~input_o ;
wire \hps_f2h_sdram0_data_writedata[223]~input_o ;
wire \hps_f2h_sdram0_data_writedata[224]~input_o ;
wire \hps_f2h_sdram0_data_writedata[225]~input_o ;
wire \hps_f2h_sdram0_data_writedata[226]~input_o ;
wire \hps_f2h_sdram0_data_writedata[227]~input_o ;
wire \hps_f2h_sdram0_data_writedata[228]~input_o ;
wire \hps_f2h_sdram0_data_writedata[229]~input_o ;
wire \hps_f2h_sdram0_data_writedata[230]~input_o ;
wire \hps_f2h_sdram0_data_writedata[231]~input_o ;
wire \hps_f2h_sdram0_data_writedata[232]~input_o ;
wire \hps_f2h_sdram0_data_writedata[233]~input_o ;
wire \hps_f2h_sdram0_data_writedata[234]~input_o ;
wire \hps_f2h_sdram0_data_writedata[235]~input_o ;
wire \hps_f2h_sdram0_data_writedata[236]~input_o ;
wire \hps_f2h_sdram0_data_writedata[237]~input_o ;
wire \hps_f2h_sdram0_data_writedata[238]~input_o ;
wire \hps_f2h_sdram0_data_writedata[239]~input_o ;
wire \hps_f2h_sdram0_data_writedata[240]~input_o ;
wire \hps_f2h_sdram0_data_writedata[241]~input_o ;
wire \hps_f2h_sdram0_data_writedata[242]~input_o ;
wire \hps_f2h_sdram0_data_writedata[243]~input_o ;
wire \hps_f2h_sdram0_data_writedata[244]~input_o ;
wire \hps_f2h_sdram0_data_writedata[245]~input_o ;
wire \hps_f2h_sdram0_data_writedata[246]~input_o ;
wire \hps_f2h_sdram0_data_writedata[247]~input_o ;
wire \hps_f2h_sdram0_data_writedata[248]~input_o ;
wire \hps_f2h_sdram0_data_writedata[249]~input_o ;
wire \hps_f2h_sdram0_data_writedata[250]~input_o ;
wire \hps_f2h_sdram0_data_writedata[251]~input_o ;
wire \hps_f2h_sdram0_data_writedata[252]~input_o ;
wire \hps_f2h_sdram0_data_writedata[253]~input_o ;
wire \hps_f2h_sdram0_data_writedata[254]~input_o ;
wire \hps_f2h_sdram0_data_writedata[255]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[24]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[25]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[26]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[27]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[28]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[29]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[30]~input_o ;
wire \hps_f2h_sdram0_data_byteenable[31]~input_o ;
wire \reset_reset_n~input_o ;
wire \state_in_export[0]~input_o ;
wire \switches_in_export[0]~input_o ;
wire \state_in_export[1]~input_o ;
wire \switches_in_export[1]~input_o ;
wire \state_in_export[2]~input_o ;
wire \switches_in_export[2]~input_o ;
wire \state_in_export[3]~input_o ;
wire \switches_in_export[3]~input_o ;
wire \state_in_export[4]~input_o ;
wire \switches_in_export[4]~input_o ;
wire \state_in_export[5]~input_o ;
wire \switches_in_export[5]~input_o ;
wire \state_in_export[6]~input_o ;
wire \switches_in_export[6]~input_o ;
wire \state_in_export[7]~input_o ;
wire \switches_in_export[7]~input_o ;
wire \state_in_export[8]~input_o ;
wire \switches_in_export[8]~input_o ;
wire \state_in_export[9]~input_o ;
wire \switches_in_export[9]~input_o ;
wire \state_in_export[10]~input_o ;
wire \state_in_export[11]~input_o ;
wire \state_in_export[12]~input_o ;
wire \state_in_export[13]~input_o ;
wire \state_in_export[14]~input_o ;
wire \state_in_export[15]~input_o ;
wire \state_in_export[16]~input_o ;
wire \state_in_export[17]~input_o ;
wire \state_in_export[18]~input_o ;
wire \state_in_export[19]~input_o ;
wire \state_in_export[20]~input_o ;
wire \state_in_export[21]~input_o ;
wire \state_in_export[22]~input_o ;
wire \state_in_export[23]~input_o ;
wire \state_in_export[24]~input_o ;
wire \state_in_export[25]~input_o ;
wire \state_in_export[26]~input_o ;
wire \state_in_export[27]~input_o ;
wire \state_in_export[28]~input_o ;
wire \state_in_export[29]~input_o ;
wire \state_in_export[30]~input_o ;
wire \state_in_export[31]~input_o ;


terminal_qsys_terminal_qsys_hps hps(
	.h2f_cold_rst_n_0(\hps|fpga_interfaces|h2f_cold_rst_n[0] ),
	.h2f_pending_rst_req_n_0(\hps|fpga_interfaces|h2f_pending_rst_req_n[0] ),
	.h2f_rst_n_0(\hps|fpga_interfaces|h2f_rst_n[0] ),
	.h2f_lw_ARVALID_0(\hps|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\hps|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\hps|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\hps|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\hps|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\hps|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\hps|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\hps|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\hps|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\hps|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\hps|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARADDR_5(\hps|fpga_interfaces|h2f_lw_ARADDR[5] ),
	.h2f_lw_ARADDR_6(\hps|fpga_interfaces|h2f_lw_ARADDR[6] ),
	.h2f_lw_ARADDR_7(\hps|fpga_interfaces|h2f_lw_ARADDR[7] ),
	.h2f_lw_ARADDR_8(\hps|fpga_interfaces|h2f_lw_ARADDR[8] ),
	.h2f_lw_ARADDR_9(\hps|fpga_interfaces|h2f_lw_ARADDR[9] ),
	.h2f_lw_ARADDR_10(\hps|fpga_interfaces|h2f_lw_ARADDR[10] ),
	.h2f_lw_ARADDR_11(\hps|fpga_interfaces|h2f_lw_ARADDR[11] ),
	.h2f_lw_ARADDR_12(\hps|fpga_interfaces|h2f_lw_ARADDR[12] ),
	.h2f_lw_ARADDR_13(\hps|fpga_interfaces|h2f_lw_ARADDR[13] ),
	.h2f_lw_ARADDR_14(\hps|fpga_interfaces|h2f_lw_ARADDR[14] ),
	.h2f_lw_ARADDR_15(\hps|fpga_interfaces|h2f_lw_ARADDR[15] ),
	.h2f_lw_ARADDR_16(\hps|fpga_interfaces|h2f_lw_ARADDR[16] ),
	.h2f_lw_ARADDR_17(\hps|fpga_interfaces|h2f_lw_ARADDR[17] ),
	.h2f_lw_ARADDR_18(\hps|fpga_interfaces|h2f_lw_ARADDR[18] ),
	.h2f_lw_ARBURST_0(\hps|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\hps|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\hps|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\hps|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\hps|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\hps|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\hps|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\hps|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\hps|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\hps|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\hps|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\hps|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\hps|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\hps|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\hps|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\hps|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\hps|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\hps|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\hps|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\hps|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\hps|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\hps|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\hps|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\hps|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\hps|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\hps|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWADDR_5(\hps|fpga_interfaces|h2f_lw_AWADDR[5] ),
	.h2f_lw_AWADDR_6(\hps|fpga_interfaces|h2f_lw_AWADDR[6] ),
	.h2f_lw_AWADDR_7(\hps|fpga_interfaces|h2f_lw_AWADDR[7] ),
	.h2f_lw_AWADDR_8(\hps|fpga_interfaces|h2f_lw_AWADDR[8] ),
	.h2f_lw_AWADDR_9(\hps|fpga_interfaces|h2f_lw_AWADDR[9] ),
	.h2f_lw_AWADDR_10(\hps|fpga_interfaces|h2f_lw_AWADDR[10] ),
	.h2f_lw_AWADDR_11(\hps|fpga_interfaces|h2f_lw_AWADDR[11] ),
	.h2f_lw_AWADDR_12(\hps|fpga_interfaces|h2f_lw_AWADDR[12] ),
	.h2f_lw_AWADDR_13(\hps|fpga_interfaces|h2f_lw_AWADDR[13] ),
	.h2f_lw_AWADDR_14(\hps|fpga_interfaces|h2f_lw_AWADDR[14] ),
	.h2f_lw_AWADDR_15(\hps|fpga_interfaces|h2f_lw_AWADDR[15] ),
	.h2f_lw_AWADDR_16(\hps|fpga_interfaces|h2f_lw_AWADDR[16] ),
	.h2f_lw_AWADDR_17(\hps|fpga_interfaces|h2f_lw_AWADDR[17] ),
	.h2f_lw_AWADDR_18(\hps|fpga_interfaces|h2f_lw_AWADDR[18] ),
	.h2f_lw_AWBURST_0(\hps|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\hps|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\hps|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\hps|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\hps|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\hps|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\hps|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\hps|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\hps|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\hps|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\hps|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\hps|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\hps|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\hps|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\hps|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\hps|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\hps|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\hps|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\hps|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\hps|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\hps|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\hps|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\hps|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\hps|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\hps|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\hps|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\hps|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\hps|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\hps|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\hps|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\hps|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\hps|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\hps|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\hps|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\hps|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\hps|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\hps|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\hps|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\hps|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\hps|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\hps|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\hps|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\hps|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\hps|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\hps|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\hps|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\hps|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\hps|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\hps|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\hps|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\hps|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\hps|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\hps|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\hps|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\hps|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\hps|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\hps|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.intermediate_1(\hps|fpga_interfaces|intermediate[1] ),
	.f2h_sdram0_READDATAVALID_0(\hps|fpga_interfaces|f2h_sdram0_READDATAVALID[0] ),
	.f2h_sdram0_READDATA_0(\hps|fpga_interfaces|f2h_sdram0_READDATA[0] ),
	.f2h_sdram0_READDATA_1(\hps|fpga_interfaces|f2h_sdram0_READDATA[1] ),
	.f2h_sdram0_READDATA_2(\hps|fpga_interfaces|f2h_sdram0_READDATA[2] ),
	.f2h_sdram0_READDATA_3(\hps|fpga_interfaces|f2h_sdram0_READDATA[3] ),
	.f2h_sdram0_READDATA_4(\hps|fpga_interfaces|f2h_sdram0_READDATA[4] ),
	.f2h_sdram0_READDATA_5(\hps|fpga_interfaces|f2h_sdram0_READDATA[5] ),
	.f2h_sdram0_READDATA_6(\hps|fpga_interfaces|f2h_sdram0_READDATA[6] ),
	.f2h_sdram0_READDATA_7(\hps|fpga_interfaces|f2h_sdram0_READDATA[7] ),
	.f2h_sdram0_READDATA_8(\hps|fpga_interfaces|f2h_sdram0_READDATA[8] ),
	.f2h_sdram0_READDATA_9(\hps|fpga_interfaces|f2h_sdram0_READDATA[9] ),
	.f2h_sdram0_READDATA_10(\hps|fpga_interfaces|f2h_sdram0_READDATA[10] ),
	.f2h_sdram0_READDATA_11(\hps|fpga_interfaces|f2h_sdram0_READDATA[11] ),
	.f2h_sdram0_READDATA_12(\hps|fpga_interfaces|f2h_sdram0_READDATA[12] ),
	.f2h_sdram0_READDATA_13(\hps|fpga_interfaces|f2h_sdram0_READDATA[13] ),
	.f2h_sdram0_READDATA_14(\hps|fpga_interfaces|f2h_sdram0_READDATA[14] ),
	.f2h_sdram0_READDATA_15(\hps|fpga_interfaces|f2h_sdram0_READDATA[15] ),
	.f2h_sdram0_READDATA_16(\hps|fpga_interfaces|f2h_sdram0_READDATA[16] ),
	.f2h_sdram0_READDATA_17(\hps|fpga_interfaces|f2h_sdram0_READDATA[17] ),
	.f2h_sdram0_READDATA_18(\hps|fpga_interfaces|f2h_sdram0_READDATA[18] ),
	.f2h_sdram0_READDATA_19(\hps|fpga_interfaces|f2h_sdram0_READDATA[19] ),
	.f2h_sdram0_READDATA_20(\hps|fpga_interfaces|f2h_sdram0_READDATA[20] ),
	.f2h_sdram0_READDATA_21(\hps|fpga_interfaces|f2h_sdram0_READDATA[21] ),
	.f2h_sdram0_READDATA_22(\hps|fpga_interfaces|f2h_sdram0_READDATA[22] ),
	.f2h_sdram0_READDATA_23(\hps|fpga_interfaces|f2h_sdram0_READDATA[23] ),
	.f2h_sdram0_READDATA_24(\hps|fpga_interfaces|f2h_sdram0_READDATA[24] ),
	.f2h_sdram0_READDATA_25(\hps|fpga_interfaces|f2h_sdram0_READDATA[25] ),
	.f2h_sdram0_READDATA_26(\hps|fpga_interfaces|f2h_sdram0_READDATA[26] ),
	.f2h_sdram0_READDATA_27(\hps|fpga_interfaces|f2h_sdram0_READDATA[27] ),
	.f2h_sdram0_READDATA_28(\hps|fpga_interfaces|f2h_sdram0_READDATA[28] ),
	.f2h_sdram0_READDATA_29(\hps|fpga_interfaces|f2h_sdram0_READDATA[29] ),
	.f2h_sdram0_READDATA_30(\hps|fpga_interfaces|f2h_sdram0_READDATA[30] ),
	.f2h_sdram0_READDATA_31(\hps|fpga_interfaces|f2h_sdram0_READDATA[31] ),
	.f2h_sdram0_READDATA_32(\hps|fpga_interfaces|f2h_sdram0_READDATA[32] ),
	.f2h_sdram0_READDATA_33(\hps|fpga_interfaces|f2h_sdram0_READDATA[33] ),
	.f2h_sdram0_READDATA_34(\hps|fpga_interfaces|f2h_sdram0_READDATA[34] ),
	.f2h_sdram0_READDATA_35(\hps|fpga_interfaces|f2h_sdram0_READDATA[35] ),
	.f2h_sdram0_READDATA_36(\hps|fpga_interfaces|f2h_sdram0_READDATA[36] ),
	.f2h_sdram0_READDATA_37(\hps|fpga_interfaces|f2h_sdram0_READDATA[37] ),
	.f2h_sdram0_READDATA_38(\hps|fpga_interfaces|f2h_sdram0_READDATA[38] ),
	.f2h_sdram0_READDATA_39(\hps|fpga_interfaces|f2h_sdram0_READDATA[39] ),
	.f2h_sdram0_READDATA_40(\hps|fpga_interfaces|f2h_sdram0_READDATA[40] ),
	.f2h_sdram0_READDATA_41(\hps|fpga_interfaces|f2h_sdram0_READDATA[41] ),
	.f2h_sdram0_READDATA_42(\hps|fpga_interfaces|f2h_sdram0_READDATA[42] ),
	.f2h_sdram0_READDATA_43(\hps|fpga_interfaces|f2h_sdram0_READDATA[43] ),
	.f2h_sdram0_READDATA_44(\hps|fpga_interfaces|f2h_sdram0_READDATA[44] ),
	.f2h_sdram0_READDATA_45(\hps|fpga_interfaces|f2h_sdram0_READDATA[45] ),
	.f2h_sdram0_READDATA_46(\hps|fpga_interfaces|f2h_sdram0_READDATA[46] ),
	.f2h_sdram0_READDATA_47(\hps|fpga_interfaces|f2h_sdram0_READDATA[47] ),
	.f2h_sdram0_READDATA_48(\hps|fpga_interfaces|f2h_sdram0_READDATA[48] ),
	.f2h_sdram0_READDATA_49(\hps|fpga_interfaces|f2h_sdram0_READDATA[49] ),
	.f2h_sdram0_READDATA_50(\hps|fpga_interfaces|f2h_sdram0_READDATA[50] ),
	.f2h_sdram0_READDATA_51(\hps|fpga_interfaces|f2h_sdram0_READDATA[51] ),
	.f2h_sdram0_READDATA_52(\hps|fpga_interfaces|f2h_sdram0_READDATA[52] ),
	.f2h_sdram0_READDATA_53(\hps|fpga_interfaces|f2h_sdram0_READDATA[53] ),
	.f2h_sdram0_READDATA_54(\hps|fpga_interfaces|f2h_sdram0_READDATA[54] ),
	.f2h_sdram0_READDATA_55(\hps|fpga_interfaces|f2h_sdram0_READDATA[55] ),
	.f2h_sdram0_READDATA_56(\hps|fpga_interfaces|f2h_sdram0_READDATA[56] ),
	.f2h_sdram0_READDATA_57(\hps|fpga_interfaces|f2h_sdram0_READDATA[57] ),
	.f2h_sdram0_READDATA_58(\hps|fpga_interfaces|f2h_sdram0_READDATA[58] ),
	.f2h_sdram0_READDATA_59(\hps|fpga_interfaces|f2h_sdram0_READDATA[59] ),
	.f2h_sdram0_READDATA_60(\hps|fpga_interfaces|f2h_sdram0_READDATA[60] ),
	.f2h_sdram0_READDATA_61(\hps|fpga_interfaces|f2h_sdram0_READDATA[61] ),
	.f2h_sdram0_READDATA_62(\hps|fpga_interfaces|f2h_sdram0_READDATA[62] ),
	.f2h_sdram0_READDATA_63(\hps|fpga_interfaces|f2h_sdram0_READDATA[63] ),
	.f2h_sdram0_READDATA_64(\hps|fpga_interfaces|f2h_sdram0_READDATA[64] ),
	.f2h_sdram0_READDATA_65(\hps|fpga_interfaces|f2h_sdram0_READDATA[65] ),
	.f2h_sdram0_READDATA_66(\hps|fpga_interfaces|f2h_sdram0_READDATA[66] ),
	.f2h_sdram0_READDATA_67(\hps|fpga_interfaces|f2h_sdram0_READDATA[67] ),
	.f2h_sdram0_READDATA_68(\hps|fpga_interfaces|f2h_sdram0_READDATA[68] ),
	.f2h_sdram0_READDATA_69(\hps|fpga_interfaces|f2h_sdram0_READDATA[69] ),
	.f2h_sdram0_READDATA_70(\hps|fpga_interfaces|f2h_sdram0_READDATA[70] ),
	.f2h_sdram0_READDATA_71(\hps|fpga_interfaces|f2h_sdram0_READDATA[71] ),
	.f2h_sdram0_READDATA_72(\hps|fpga_interfaces|f2h_sdram0_READDATA[72] ),
	.f2h_sdram0_READDATA_73(\hps|fpga_interfaces|f2h_sdram0_READDATA[73] ),
	.f2h_sdram0_READDATA_74(\hps|fpga_interfaces|f2h_sdram0_READDATA[74] ),
	.f2h_sdram0_READDATA_75(\hps|fpga_interfaces|f2h_sdram0_READDATA[75] ),
	.f2h_sdram0_READDATA_76(\hps|fpga_interfaces|f2h_sdram0_READDATA[76] ),
	.f2h_sdram0_READDATA_77(\hps|fpga_interfaces|f2h_sdram0_READDATA[77] ),
	.f2h_sdram0_READDATA_78(\hps|fpga_interfaces|f2h_sdram0_READDATA[78] ),
	.f2h_sdram0_READDATA_79(\hps|fpga_interfaces|f2h_sdram0_READDATA[79] ),
	.f2h_sdram0_READDATA_80(\hps|fpga_interfaces|f2h_sdram0_READDATA[80] ),
	.f2h_sdram0_READDATA_81(\hps|fpga_interfaces|f2h_sdram0_READDATA[81] ),
	.f2h_sdram0_READDATA_82(\hps|fpga_interfaces|f2h_sdram0_READDATA[82] ),
	.f2h_sdram0_READDATA_83(\hps|fpga_interfaces|f2h_sdram0_READDATA[83] ),
	.f2h_sdram0_READDATA_84(\hps|fpga_interfaces|f2h_sdram0_READDATA[84] ),
	.f2h_sdram0_READDATA_85(\hps|fpga_interfaces|f2h_sdram0_READDATA[85] ),
	.f2h_sdram0_READDATA_86(\hps|fpga_interfaces|f2h_sdram0_READDATA[86] ),
	.f2h_sdram0_READDATA_87(\hps|fpga_interfaces|f2h_sdram0_READDATA[87] ),
	.f2h_sdram0_READDATA_88(\hps|fpga_interfaces|f2h_sdram0_READDATA[88] ),
	.f2h_sdram0_READDATA_89(\hps|fpga_interfaces|f2h_sdram0_READDATA[89] ),
	.f2h_sdram0_READDATA_90(\hps|fpga_interfaces|f2h_sdram0_READDATA[90] ),
	.f2h_sdram0_READDATA_91(\hps|fpga_interfaces|f2h_sdram0_READDATA[91] ),
	.f2h_sdram0_READDATA_92(\hps|fpga_interfaces|f2h_sdram0_READDATA[92] ),
	.f2h_sdram0_READDATA_93(\hps|fpga_interfaces|f2h_sdram0_READDATA[93] ),
	.f2h_sdram0_READDATA_94(\hps|fpga_interfaces|f2h_sdram0_READDATA[94] ),
	.f2h_sdram0_READDATA_95(\hps|fpga_interfaces|f2h_sdram0_READDATA[95] ),
	.f2h_sdram0_READDATA_96(\hps|fpga_interfaces|f2h_sdram0_READDATA[96] ),
	.f2h_sdram0_READDATA_97(\hps|fpga_interfaces|f2h_sdram0_READDATA[97] ),
	.f2h_sdram0_READDATA_98(\hps|fpga_interfaces|f2h_sdram0_READDATA[98] ),
	.f2h_sdram0_READDATA_99(\hps|fpga_interfaces|f2h_sdram0_READDATA[99] ),
	.f2h_sdram0_READDATA_100(\hps|fpga_interfaces|f2h_sdram0_READDATA[100] ),
	.f2h_sdram0_READDATA_101(\hps|fpga_interfaces|f2h_sdram0_READDATA[101] ),
	.f2h_sdram0_READDATA_102(\hps|fpga_interfaces|f2h_sdram0_READDATA[102] ),
	.f2h_sdram0_READDATA_103(\hps|fpga_interfaces|f2h_sdram0_READDATA[103] ),
	.f2h_sdram0_READDATA_104(\hps|fpga_interfaces|f2h_sdram0_READDATA[104] ),
	.f2h_sdram0_READDATA_105(\hps|fpga_interfaces|f2h_sdram0_READDATA[105] ),
	.f2h_sdram0_READDATA_106(\hps|fpga_interfaces|f2h_sdram0_READDATA[106] ),
	.f2h_sdram0_READDATA_107(\hps|fpga_interfaces|f2h_sdram0_READDATA[107] ),
	.f2h_sdram0_READDATA_108(\hps|fpga_interfaces|f2h_sdram0_READDATA[108] ),
	.f2h_sdram0_READDATA_109(\hps|fpga_interfaces|f2h_sdram0_READDATA[109] ),
	.f2h_sdram0_READDATA_110(\hps|fpga_interfaces|f2h_sdram0_READDATA[110] ),
	.f2h_sdram0_READDATA_111(\hps|fpga_interfaces|f2h_sdram0_READDATA[111] ),
	.f2h_sdram0_READDATA_112(\hps|fpga_interfaces|f2h_sdram0_READDATA[112] ),
	.f2h_sdram0_READDATA_113(\hps|fpga_interfaces|f2h_sdram0_READDATA[113] ),
	.f2h_sdram0_READDATA_114(\hps|fpga_interfaces|f2h_sdram0_READDATA[114] ),
	.f2h_sdram0_READDATA_115(\hps|fpga_interfaces|f2h_sdram0_READDATA[115] ),
	.f2h_sdram0_READDATA_116(\hps|fpga_interfaces|f2h_sdram0_READDATA[116] ),
	.f2h_sdram0_READDATA_117(\hps|fpga_interfaces|f2h_sdram0_READDATA[117] ),
	.f2h_sdram0_READDATA_118(\hps|fpga_interfaces|f2h_sdram0_READDATA[118] ),
	.f2h_sdram0_READDATA_119(\hps|fpga_interfaces|f2h_sdram0_READDATA[119] ),
	.f2h_sdram0_READDATA_120(\hps|fpga_interfaces|f2h_sdram0_READDATA[120] ),
	.f2h_sdram0_READDATA_121(\hps|fpga_interfaces|f2h_sdram0_READDATA[121] ),
	.f2h_sdram0_READDATA_122(\hps|fpga_interfaces|f2h_sdram0_READDATA[122] ),
	.f2h_sdram0_READDATA_123(\hps|fpga_interfaces|f2h_sdram0_READDATA[123] ),
	.f2h_sdram0_READDATA_124(\hps|fpga_interfaces|f2h_sdram0_READDATA[124] ),
	.f2h_sdram0_READDATA_125(\hps|fpga_interfaces|f2h_sdram0_READDATA[125] ),
	.f2h_sdram0_READDATA_126(\hps|fpga_interfaces|f2h_sdram0_READDATA[126] ),
	.f2h_sdram0_READDATA_127(\hps|fpga_interfaces|f2h_sdram0_READDATA[127] ),
	.f2h_sdram0_READDATA_128(\hps|fpga_interfaces|f2h_sdram0_READDATA[128] ),
	.f2h_sdram0_READDATA_129(\hps|fpga_interfaces|f2h_sdram0_READDATA[129] ),
	.f2h_sdram0_READDATA_130(\hps|fpga_interfaces|f2h_sdram0_READDATA[130] ),
	.f2h_sdram0_READDATA_131(\hps|fpga_interfaces|f2h_sdram0_READDATA[131] ),
	.f2h_sdram0_READDATA_132(\hps|fpga_interfaces|f2h_sdram0_READDATA[132] ),
	.f2h_sdram0_READDATA_133(\hps|fpga_interfaces|f2h_sdram0_READDATA[133] ),
	.f2h_sdram0_READDATA_134(\hps|fpga_interfaces|f2h_sdram0_READDATA[134] ),
	.f2h_sdram0_READDATA_135(\hps|fpga_interfaces|f2h_sdram0_READDATA[135] ),
	.f2h_sdram0_READDATA_136(\hps|fpga_interfaces|f2h_sdram0_READDATA[136] ),
	.f2h_sdram0_READDATA_137(\hps|fpga_interfaces|f2h_sdram0_READDATA[137] ),
	.f2h_sdram0_READDATA_138(\hps|fpga_interfaces|f2h_sdram0_READDATA[138] ),
	.f2h_sdram0_READDATA_139(\hps|fpga_interfaces|f2h_sdram0_READDATA[139] ),
	.f2h_sdram0_READDATA_140(\hps|fpga_interfaces|f2h_sdram0_READDATA[140] ),
	.f2h_sdram0_READDATA_141(\hps|fpga_interfaces|f2h_sdram0_READDATA[141] ),
	.f2h_sdram0_READDATA_142(\hps|fpga_interfaces|f2h_sdram0_READDATA[142] ),
	.f2h_sdram0_READDATA_143(\hps|fpga_interfaces|f2h_sdram0_READDATA[143] ),
	.f2h_sdram0_READDATA_144(\hps|fpga_interfaces|f2h_sdram0_READDATA[144] ),
	.f2h_sdram0_READDATA_145(\hps|fpga_interfaces|f2h_sdram0_READDATA[145] ),
	.f2h_sdram0_READDATA_146(\hps|fpga_interfaces|f2h_sdram0_READDATA[146] ),
	.f2h_sdram0_READDATA_147(\hps|fpga_interfaces|f2h_sdram0_READDATA[147] ),
	.f2h_sdram0_READDATA_148(\hps|fpga_interfaces|f2h_sdram0_READDATA[148] ),
	.f2h_sdram0_READDATA_149(\hps|fpga_interfaces|f2h_sdram0_READDATA[149] ),
	.f2h_sdram0_READDATA_150(\hps|fpga_interfaces|f2h_sdram0_READDATA[150] ),
	.f2h_sdram0_READDATA_151(\hps|fpga_interfaces|f2h_sdram0_READDATA[151] ),
	.f2h_sdram0_READDATA_152(\hps|fpga_interfaces|f2h_sdram0_READDATA[152] ),
	.f2h_sdram0_READDATA_153(\hps|fpga_interfaces|f2h_sdram0_READDATA[153] ),
	.f2h_sdram0_READDATA_154(\hps|fpga_interfaces|f2h_sdram0_READDATA[154] ),
	.f2h_sdram0_READDATA_155(\hps|fpga_interfaces|f2h_sdram0_READDATA[155] ),
	.f2h_sdram0_READDATA_156(\hps|fpga_interfaces|f2h_sdram0_READDATA[156] ),
	.f2h_sdram0_READDATA_157(\hps|fpga_interfaces|f2h_sdram0_READDATA[157] ),
	.f2h_sdram0_READDATA_158(\hps|fpga_interfaces|f2h_sdram0_READDATA[158] ),
	.f2h_sdram0_READDATA_159(\hps|fpga_interfaces|f2h_sdram0_READDATA[159] ),
	.f2h_sdram0_READDATA_160(\hps|fpga_interfaces|f2h_sdram0_READDATA[160] ),
	.f2h_sdram0_READDATA_161(\hps|fpga_interfaces|f2h_sdram0_READDATA[161] ),
	.f2h_sdram0_READDATA_162(\hps|fpga_interfaces|f2h_sdram0_READDATA[162] ),
	.f2h_sdram0_READDATA_163(\hps|fpga_interfaces|f2h_sdram0_READDATA[163] ),
	.f2h_sdram0_READDATA_164(\hps|fpga_interfaces|f2h_sdram0_READDATA[164] ),
	.f2h_sdram0_READDATA_165(\hps|fpga_interfaces|f2h_sdram0_READDATA[165] ),
	.f2h_sdram0_READDATA_166(\hps|fpga_interfaces|f2h_sdram0_READDATA[166] ),
	.f2h_sdram0_READDATA_167(\hps|fpga_interfaces|f2h_sdram0_READDATA[167] ),
	.f2h_sdram0_READDATA_168(\hps|fpga_interfaces|f2h_sdram0_READDATA[168] ),
	.f2h_sdram0_READDATA_169(\hps|fpga_interfaces|f2h_sdram0_READDATA[169] ),
	.f2h_sdram0_READDATA_170(\hps|fpga_interfaces|f2h_sdram0_READDATA[170] ),
	.f2h_sdram0_READDATA_171(\hps|fpga_interfaces|f2h_sdram0_READDATA[171] ),
	.f2h_sdram0_READDATA_172(\hps|fpga_interfaces|f2h_sdram0_READDATA[172] ),
	.f2h_sdram0_READDATA_173(\hps|fpga_interfaces|f2h_sdram0_READDATA[173] ),
	.f2h_sdram0_READDATA_174(\hps|fpga_interfaces|f2h_sdram0_READDATA[174] ),
	.f2h_sdram0_READDATA_175(\hps|fpga_interfaces|f2h_sdram0_READDATA[175] ),
	.f2h_sdram0_READDATA_176(\hps|fpga_interfaces|f2h_sdram0_READDATA[176] ),
	.f2h_sdram0_READDATA_177(\hps|fpga_interfaces|f2h_sdram0_READDATA[177] ),
	.f2h_sdram0_READDATA_178(\hps|fpga_interfaces|f2h_sdram0_READDATA[178] ),
	.f2h_sdram0_READDATA_179(\hps|fpga_interfaces|f2h_sdram0_READDATA[179] ),
	.f2h_sdram0_READDATA_180(\hps|fpga_interfaces|f2h_sdram0_READDATA[180] ),
	.f2h_sdram0_READDATA_181(\hps|fpga_interfaces|f2h_sdram0_READDATA[181] ),
	.f2h_sdram0_READDATA_182(\hps|fpga_interfaces|f2h_sdram0_READDATA[182] ),
	.f2h_sdram0_READDATA_183(\hps|fpga_interfaces|f2h_sdram0_READDATA[183] ),
	.f2h_sdram0_READDATA_184(\hps|fpga_interfaces|f2h_sdram0_READDATA[184] ),
	.f2h_sdram0_READDATA_185(\hps|fpga_interfaces|f2h_sdram0_READDATA[185] ),
	.f2h_sdram0_READDATA_186(\hps|fpga_interfaces|f2h_sdram0_READDATA[186] ),
	.f2h_sdram0_READDATA_187(\hps|fpga_interfaces|f2h_sdram0_READDATA[187] ),
	.f2h_sdram0_READDATA_188(\hps|fpga_interfaces|f2h_sdram0_READDATA[188] ),
	.f2h_sdram0_READDATA_189(\hps|fpga_interfaces|f2h_sdram0_READDATA[189] ),
	.f2h_sdram0_READDATA_190(\hps|fpga_interfaces|f2h_sdram0_READDATA[190] ),
	.f2h_sdram0_READDATA_191(\hps|fpga_interfaces|f2h_sdram0_READDATA[191] ),
	.f2h_sdram0_READDATA_192(\hps|fpga_interfaces|f2h_sdram0_READDATA[192] ),
	.f2h_sdram0_READDATA_193(\hps|fpga_interfaces|f2h_sdram0_READDATA[193] ),
	.f2h_sdram0_READDATA_194(\hps|fpga_interfaces|f2h_sdram0_READDATA[194] ),
	.f2h_sdram0_READDATA_195(\hps|fpga_interfaces|f2h_sdram0_READDATA[195] ),
	.f2h_sdram0_READDATA_196(\hps|fpga_interfaces|f2h_sdram0_READDATA[196] ),
	.f2h_sdram0_READDATA_197(\hps|fpga_interfaces|f2h_sdram0_READDATA[197] ),
	.f2h_sdram0_READDATA_198(\hps|fpga_interfaces|f2h_sdram0_READDATA[198] ),
	.f2h_sdram0_READDATA_199(\hps|fpga_interfaces|f2h_sdram0_READDATA[199] ),
	.f2h_sdram0_READDATA_200(\hps|fpga_interfaces|f2h_sdram0_READDATA[200] ),
	.f2h_sdram0_READDATA_201(\hps|fpga_interfaces|f2h_sdram0_READDATA[201] ),
	.f2h_sdram0_READDATA_202(\hps|fpga_interfaces|f2h_sdram0_READDATA[202] ),
	.f2h_sdram0_READDATA_203(\hps|fpga_interfaces|f2h_sdram0_READDATA[203] ),
	.f2h_sdram0_READDATA_204(\hps|fpga_interfaces|f2h_sdram0_READDATA[204] ),
	.f2h_sdram0_READDATA_205(\hps|fpga_interfaces|f2h_sdram0_READDATA[205] ),
	.f2h_sdram0_READDATA_206(\hps|fpga_interfaces|f2h_sdram0_READDATA[206] ),
	.f2h_sdram0_READDATA_207(\hps|fpga_interfaces|f2h_sdram0_READDATA[207] ),
	.f2h_sdram0_READDATA_208(\hps|fpga_interfaces|f2h_sdram0_READDATA[208] ),
	.f2h_sdram0_READDATA_209(\hps|fpga_interfaces|f2h_sdram0_READDATA[209] ),
	.f2h_sdram0_READDATA_210(\hps|fpga_interfaces|f2h_sdram0_READDATA[210] ),
	.f2h_sdram0_READDATA_211(\hps|fpga_interfaces|f2h_sdram0_READDATA[211] ),
	.f2h_sdram0_READDATA_212(\hps|fpga_interfaces|f2h_sdram0_READDATA[212] ),
	.f2h_sdram0_READDATA_213(\hps|fpga_interfaces|f2h_sdram0_READDATA[213] ),
	.f2h_sdram0_READDATA_214(\hps|fpga_interfaces|f2h_sdram0_READDATA[214] ),
	.f2h_sdram0_READDATA_215(\hps|fpga_interfaces|f2h_sdram0_READDATA[215] ),
	.f2h_sdram0_READDATA_216(\hps|fpga_interfaces|f2h_sdram0_READDATA[216] ),
	.f2h_sdram0_READDATA_217(\hps|fpga_interfaces|f2h_sdram0_READDATA[217] ),
	.f2h_sdram0_READDATA_218(\hps|fpga_interfaces|f2h_sdram0_READDATA[218] ),
	.f2h_sdram0_READDATA_219(\hps|fpga_interfaces|f2h_sdram0_READDATA[219] ),
	.f2h_sdram0_READDATA_220(\hps|fpga_interfaces|f2h_sdram0_READDATA[220] ),
	.f2h_sdram0_READDATA_221(\hps|fpga_interfaces|f2h_sdram0_READDATA[221] ),
	.f2h_sdram0_READDATA_222(\hps|fpga_interfaces|f2h_sdram0_READDATA[222] ),
	.f2h_sdram0_READDATA_223(\hps|fpga_interfaces|f2h_sdram0_READDATA[223] ),
	.f2h_sdram0_READDATA_224(\hps|fpga_interfaces|f2h_sdram0_READDATA[224] ),
	.f2h_sdram0_READDATA_225(\hps|fpga_interfaces|f2h_sdram0_READDATA[225] ),
	.f2h_sdram0_READDATA_226(\hps|fpga_interfaces|f2h_sdram0_READDATA[226] ),
	.f2h_sdram0_READDATA_227(\hps|fpga_interfaces|f2h_sdram0_READDATA[227] ),
	.f2h_sdram0_READDATA_228(\hps|fpga_interfaces|f2h_sdram0_READDATA[228] ),
	.f2h_sdram0_READDATA_229(\hps|fpga_interfaces|f2h_sdram0_READDATA[229] ),
	.f2h_sdram0_READDATA_230(\hps|fpga_interfaces|f2h_sdram0_READDATA[230] ),
	.f2h_sdram0_READDATA_231(\hps|fpga_interfaces|f2h_sdram0_READDATA[231] ),
	.f2h_sdram0_READDATA_232(\hps|fpga_interfaces|f2h_sdram0_READDATA[232] ),
	.f2h_sdram0_READDATA_233(\hps|fpga_interfaces|f2h_sdram0_READDATA[233] ),
	.f2h_sdram0_READDATA_234(\hps|fpga_interfaces|f2h_sdram0_READDATA[234] ),
	.f2h_sdram0_READDATA_235(\hps|fpga_interfaces|f2h_sdram0_READDATA[235] ),
	.f2h_sdram0_READDATA_236(\hps|fpga_interfaces|f2h_sdram0_READDATA[236] ),
	.f2h_sdram0_READDATA_237(\hps|fpga_interfaces|f2h_sdram0_READDATA[237] ),
	.f2h_sdram0_READDATA_238(\hps|fpga_interfaces|f2h_sdram0_READDATA[238] ),
	.f2h_sdram0_READDATA_239(\hps|fpga_interfaces|f2h_sdram0_READDATA[239] ),
	.f2h_sdram0_READDATA_240(\hps|fpga_interfaces|f2h_sdram0_READDATA[240] ),
	.f2h_sdram0_READDATA_241(\hps|fpga_interfaces|f2h_sdram0_READDATA[241] ),
	.f2h_sdram0_READDATA_242(\hps|fpga_interfaces|f2h_sdram0_READDATA[242] ),
	.f2h_sdram0_READDATA_243(\hps|fpga_interfaces|f2h_sdram0_READDATA[243] ),
	.f2h_sdram0_READDATA_244(\hps|fpga_interfaces|f2h_sdram0_READDATA[244] ),
	.f2h_sdram0_READDATA_245(\hps|fpga_interfaces|f2h_sdram0_READDATA[245] ),
	.f2h_sdram0_READDATA_246(\hps|fpga_interfaces|f2h_sdram0_READDATA[246] ),
	.f2h_sdram0_READDATA_247(\hps|fpga_interfaces|f2h_sdram0_READDATA[247] ),
	.f2h_sdram0_READDATA_248(\hps|fpga_interfaces|f2h_sdram0_READDATA[248] ),
	.f2h_sdram0_READDATA_249(\hps|fpga_interfaces|f2h_sdram0_READDATA[249] ),
	.f2h_sdram0_READDATA_250(\hps|fpga_interfaces|f2h_sdram0_READDATA[250] ),
	.f2h_sdram0_READDATA_251(\hps|fpga_interfaces|f2h_sdram0_READDATA[251] ),
	.f2h_sdram0_READDATA_252(\hps|fpga_interfaces|f2h_sdram0_READDATA[252] ),
	.f2h_sdram0_READDATA_253(\hps|fpga_interfaces|f2h_sdram0_READDATA[253] ),
	.f2h_sdram0_READDATA_254(\hps|fpga_interfaces|f2h_sdram0_READDATA[254] ),
	.f2h_sdram0_READDATA_255(\hps|fpga_interfaces|f2h_sdram0_READDATA[255] ),
	.cmd_sink_ready(\mm_interconnect_0|hps_h2f_lw_axi_master_rd_limiter|cmd_sink_ready~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.nonposted_cmd_accepted1(\mm_interconnect_0|hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~5_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux_001|src_data[1]~11_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~17_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux_001|src_data[3]~23_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux_001|src_data[4]~29_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~35_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~41_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~48_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~54_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~58_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux_001|src_payload~11_combout ),
	.src_payload13(\mm_interconnect_0|rsp_mux_001|src_payload~14_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux_001|src_payload~17_combout ),
	.src_payload15(\mm_interconnect_0|rsp_mux_001|src_payload~20_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux_001|src_payload~23_combout ),
	.src_payload17(\mm_interconnect_0|rsp_mux_001|src_payload~26_combout ),
	.src_payload18(\mm_interconnect_0|rsp_mux_001|src_payload~29_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux_001|src_payload~32_combout ),
	.src_payload20(\mm_interconnect_0|rsp_mux_001|src_payload~35_combout ),
	.src_payload21(\mm_interconnect_0|rsp_mux_001|src_payload~38_combout ),
	.src_payload22(\mm_interconnect_0|rsp_mux_001|src_payload~41_combout ),
	.src_payload23(\mm_interconnect_0|rsp_mux_001|src_payload~44_combout ),
	.src_payload24(\mm_interconnect_0|rsp_mux_001|src_payload~47_combout ),
	.src_payload25(\mm_interconnect_0|rsp_mux_001|src_payload~50_combout ),
	.src_payload26(\mm_interconnect_0|rsp_mux_001|src_payload~53_combout ),
	.src_payload27(\mm_interconnect_0|rsp_mux_001|src_payload~56_combout ),
	.src_payload28(\mm_interconnect_0|rsp_mux_001|src_payload~59_combout ),
	.src_payload29(\mm_interconnect_0|rsp_mux_001|src_payload~62_combout ),
	.src_payload30(\mm_interconnect_0|rsp_mux_001|src_payload~65_combout ),
	.src_payload31(\mm_interconnect_0|rsp_mux_001|src_payload~68_combout ),
	.src_payload32(\mm_interconnect_0|rsp_mux_001|src_payload~71_combout ),
	.src_payload33(\mm_interconnect_0|rsp_mux_001|src_payload~74_combout ),
	.src_data_92(\mm_interconnect_0|rsp_mux_001|src_data[92]~combout ),
	.src_data_93(\mm_interconnect_0|rsp_mux_001|src_data[93]~combout ),
	.src_data_94(\mm_interconnect_0|rsp_mux_001|src_data[94]~combout ),
	.src_data_95(\mm_interconnect_0|rsp_mux_001|src_data[95]~combout ),
	.src_data_96(\mm_interconnect_0|rsp_mux_001|src_data[96]~combout ),
	.src_data_97(\mm_interconnect_0|rsp_mux_001|src_data[97]~combout ),
	.src_data_98(\mm_interconnect_0|rsp_mux_001|src_data[98]~combout ),
	.src_data_99(\mm_interconnect_0|rsp_mux_001|src_data[99]~combout ),
	.src_data_100(\mm_interconnect_0|rsp_mux_001|src_data[100]~combout ),
	.src_data_101(\mm_interconnect_0|rsp_mux_001|src_data[101]~combout ),
	.src_data_102(\mm_interconnect_0|rsp_mux_001|src_data[102]~combout ),
	.src_data_103(\mm_interconnect_0|rsp_mux_001|src_data[103]~combout ),
	.emac1_inst(\hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ),
	.emac1_inst1(\hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ),
	.intermediate_0(\hps|hps_io|border|intermediate[0] ),
	.intermediate_11(\hps|hps_io|border|intermediate[1] ),
	.emac1_inst2(\hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ),
	.emac1_inst3(\hps|hps_io|border|emac1_inst~emac_phy_txd ),
	.emac1_inst4(\hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ),
	.emac1_inst5(\hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ),
	.emac1_inst6(\hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ),
	.sdio_inst(\hps|hps_io|border|sdio_inst~sdmmc_cclk ),
	.intermediate_2(\hps|hps_io|border|intermediate[2] ),
	.intermediate_3(\hps|hps_io|border|intermediate[3] ),
	.intermediate_4(\hps|hps_io|border|intermediate[4] ),
	.intermediate_6(\hps|hps_io|border|intermediate[6] ),
	.intermediate_8(\hps|hps_io|border|intermediate[8] ),
	.intermediate_10(\hps|hps_io|border|intermediate[10] ),
	.intermediate_5(\hps|hps_io|border|intermediate[5] ),
	.intermediate_7(\hps|hps_io|border|intermediate[7] ),
	.intermediate_9(\hps|hps_io|border|intermediate[9] ),
	.intermediate_111(\hps|hps_io|border|intermediate[11] ),
	.uart0_inst(\hps|hps_io|border|uart0_inst~uart_txd ),
	.parallelterminationcontrol_0(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] ),
	.parallelterminationcontrol_1(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ),
	.parallelterminationcontrol_2(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ),
	.parallelterminationcontrol_3(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ),
	.parallelterminationcontrol_4(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ),
	.parallelterminationcontrol_5(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ),
	.parallelterminationcontrol_6(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ),
	.parallelterminationcontrol_7(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ),
	.parallelterminationcontrol_8(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ),
	.parallelterminationcontrol_9(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ),
	.parallelterminationcontrol_10(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ),
	.parallelterminationcontrol_11(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ),
	.parallelterminationcontrol_12(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ),
	.parallelterminationcontrol_13(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ),
	.parallelterminationcontrol_14(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ),
	.parallelterminationcontrol_15(\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ),
	.seriesterminationcontrol_0(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] ),
	.seriesterminationcontrol_1(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ),
	.seriesterminationcontrol_2(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ),
	.seriesterminationcontrol_3(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ),
	.seriesterminationcontrol_4(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ),
	.seriesterminationcontrol_5(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ),
	.seriesterminationcontrol_6(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ),
	.seriesterminationcontrol_7(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ),
	.seriesterminationcontrol_8(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ),
	.seriesterminationcontrol_9(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ),
	.seriesterminationcontrol_10(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ),
	.seriesterminationcontrol_11(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ),
	.seriesterminationcontrol_12(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ),
	.seriesterminationcontrol_13(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ),
	.seriesterminationcontrol_14(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ),
	.seriesterminationcontrol_15(\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ),
	.dqsin(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dqsin3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ),
	.pad_gen0raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ),
	.pad_gen1raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ),
	.pad_gen2raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ),
	.pad_gen3raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ),
	.pad_gen4raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ),
	.pad_gen5raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ),
	.pad_gen6raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ),
	.pad_gen7raw_input3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ),
	.dataout_0(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ),
	.dataout_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ),
	.dataout_2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ),
	.dataout_3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ),
	.dataout_4(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ),
	.dataout_5(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ),
	.dataout_6(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ),
	.dataout_7(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ),
	.dataout_8(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ),
	.dataout_9(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ),
	.dataout_10(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ),
	.dataout_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ),
	.dataout_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ),
	.dataout_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ),
	.dataout_14(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ),
	.dataout_01(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ),
	.dataout_15(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ),
	.dataout_21(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ),
	.dataout_16(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ),
	.dataout_02(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ),
	.dataout_31(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ),
	.dataout_41(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ),
	.dataout_51(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ),
	.dataout_03(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ),
	.dataout_22(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ),
	.extra_output_pad_gen0delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.extra_output_pad_gen0delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.wire_pseudo_diffa_o_0(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.wire_pseudo_diffa_obar_0(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.wire_pseudo_diffa_oeout_0(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.wire_pseudo_diffa_oebout_0(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.pad_gen0delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_11(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_12(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.pad_gen0delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.pad_gen0delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.delayed_oct3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.pad_gen1delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.pad_gen1delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.pad_gen2delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.pad_gen2delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.pad_gen3delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.pad_gen3delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.pad_gen4delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.pad_gen4delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.pad_gen5delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.pad_gen5delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.pad_gen6delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.pad_gen6delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.pad_gen7delayed_data_out3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.pad_gen7delayed_oe_13(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.os(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar1(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar2(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.os3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.os_bar3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.diff_oe3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.diff_oe_bar3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.diff_dtc3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.diff_dtc_bar3(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.hps_io_emac1_inst_MDIO_0(\hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o ),
	.hps_io_sdio_inst_CMD_0(\hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o ),
	.hps_io_sdio_inst_D0_0(\hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o ),
	.hps_io_sdio_inst_D1_0(\hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o ),
	.hps_io_sdio_inst_D2_0(\hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o ),
	.hps_io_sdio_inst_D3_0(\hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_0(\hps_f2h_stm_hw_events_stm_hwevents[0]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_1(\hps_f2h_stm_hw_events_stm_hwevents[1]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_2(\hps_f2h_stm_hw_events_stm_hwevents[2]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_3(\hps_f2h_stm_hw_events_stm_hwevents[3]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_4(\hps_f2h_stm_hw_events_stm_hwevents[4]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_5(\hps_f2h_stm_hw_events_stm_hwevents[5]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_6(\hps_f2h_stm_hw_events_stm_hwevents[6]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_7(\hps_f2h_stm_hw_events_stm_hwevents[7]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_8(\hps_f2h_stm_hw_events_stm_hwevents[8]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_9(\hps_f2h_stm_hw_events_stm_hwevents[9]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_10(\hps_f2h_stm_hw_events_stm_hwevents[10]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_11(\hps_f2h_stm_hw_events_stm_hwevents[11]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_12(\hps_f2h_stm_hw_events_stm_hwevents[12]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_13(\hps_f2h_stm_hw_events_stm_hwevents[13]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_14(\hps_f2h_stm_hw_events_stm_hwevents[14]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_15(\hps_f2h_stm_hw_events_stm_hwevents[15]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_16(\hps_f2h_stm_hw_events_stm_hwevents[16]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_17(\hps_f2h_stm_hw_events_stm_hwevents[17]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_18(\hps_f2h_stm_hw_events_stm_hwevents[18]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_19(\hps_f2h_stm_hw_events_stm_hwevents[19]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_20(\hps_f2h_stm_hw_events_stm_hwevents[20]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_21(\hps_f2h_stm_hw_events_stm_hwevents[21]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_22(\hps_f2h_stm_hw_events_stm_hwevents[22]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_23(\hps_f2h_stm_hw_events_stm_hwevents[23]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_24(\hps_f2h_stm_hw_events_stm_hwevents[24]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_25(\hps_f2h_stm_hw_events_stm_hwevents[25]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_26(\hps_f2h_stm_hw_events_stm_hwevents[26]~input_o ),
	.hps_f2h_stm_hw_events_stm_hwevents_27(\hps_f2h_stm_hw_events_stm_hwevents[27]~input_o ),
	.clk_clk(\clk_clk~input_o ),
	.hps_hps_io_hps_io_emac1_inst_RXD0(\hps_hps_io_hps_io_emac1_inst_RXD0~input_o ),
	.hps_hps_io_hps_io_emac1_inst_RXD1(\hps_hps_io_hps_io_emac1_inst_RXD1~input_o ),
	.hps_hps_io_hps_io_emac1_inst_RXD2(\hps_hps_io_hps_io_emac1_inst_RXD2~input_o ),
	.hps_hps_io_hps_io_emac1_inst_RXD3(\hps_hps_io_hps_io_emac1_inst_RXD3~input_o ),
	.hps_hps_io_hps_io_emac1_inst_RX_CLK(\hps_hps_io_hps_io_emac1_inst_RX_CLK~input_o ),
	.hps_hps_io_hps_io_emac1_inst_RX_CTL(\hps_hps_io_hps_io_emac1_inst_RX_CTL~input_o ),
	.hps_hps_io_hps_io_uart0_inst_RX(\hps_hps_io_hps_io_uart0_inst_RX~input_o ),
	.memory_oct_rzqin(\memory_oct_rzqin~input_o ),
	.hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n(\hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n~input_o ),
	.hps_f2h_sdram0_data_read(\hps_f2h_sdram0_data_read~input_o ),
	.hps_f2h_sdram0_data_write(\hps_f2h_sdram0_data_write~input_o ),
	.hps_f2h_sdram0_data_address_0(\hps_f2h_sdram0_data_address[0]~input_o ),
	.hps_f2h_sdram0_data_address_1(\hps_f2h_sdram0_data_address[1]~input_o ),
	.hps_f2h_sdram0_data_address_2(\hps_f2h_sdram0_data_address[2]~input_o ),
	.hps_f2h_sdram0_data_address_3(\hps_f2h_sdram0_data_address[3]~input_o ),
	.hps_f2h_sdram0_data_address_4(\hps_f2h_sdram0_data_address[4]~input_o ),
	.hps_f2h_sdram0_data_address_5(\hps_f2h_sdram0_data_address[5]~input_o ),
	.hps_f2h_sdram0_data_address_6(\hps_f2h_sdram0_data_address[6]~input_o ),
	.hps_f2h_sdram0_data_address_7(\hps_f2h_sdram0_data_address[7]~input_o ),
	.hps_f2h_sdram0_data_address_8(\hps_f2h_sdram0_data_address[8]~input_o ),
	.hps_f2h_sdram0_data_address_9(\hps_f2h_sdram0_data_address[9]~input_o ),
	.hps_f2h_sdram0_data_address_10(\hps_f2h_sdram0_data_address[10]~input_o ),
	.hps_f2h_sdram0_data_address_11(\hps_f2h_sdram0_data_address[11]~input_o ),
	.hps_f2h_sdram0_data_address_12(\hps_f2h_sdram0_data_address[12]~input_o ),
	.hps_f2h_sdram0_data_address_13(\hps_f2h_sdram0_data_address[13]~input_o ),
	.hps_f2h_sdram0_data_address_14(\hps_f2h_sdram0_data_address[14]~input_o ),
	.hps_f2h_sdram0_data_address_15(\hps_f2h_sdram0_data_address[15]~input_o ),
	.hps_f2h_sdram0_data_address_16(\hps_f2h_sdram0_data_address[16]~input_o ),
	.hps_f2h_sdram0_data_address_17(\hps_f2h_sdram0_data_address[17]~input_o ),
	.hps_f2h_sdram0_data_address_18(\hps_f2h_sdram0_data_address[18]~input_o ),
	.hps_f2h_sdram0_data_address_19(\hps_f2h_sdram0_data_address[19]~input_o ),
	.hps_f2h_sdram0_data_address_20(\hps_f2h_sdram0_data_address[20]~input_o ),
	.hps_f2h_sdram0_data_address_21(\hps_f2h_sdram0_data_address[21]~input_o ),
	.hps_f2h_sdram0_data_address_22(\hps_f2h_sdram0_data_address[22]~input_o ),
	.hps_f2h_sdram0_data_address_23(\hps_f2h_sdram0_data_address[23]~input_o ),
	.hps_f2h_sdram0_data_address_24(\hps_f2h_sdram0_data_address[24]~input_o ),
	.hps_f2h_sdram0_data_address_25(\hps_f2h_sdram0_data_address[25]~input_o ),
	.hps_f2h_sdram0_data_address_26(\hps_f2h_sdram0_data_address[26]~input_o ),
	.hps_f2h_sdram0_data_burstcount_0(\hps_f2h_sdram0_data_burstcount[0]~input_o ),
	.hps_f2h_sdram0_data_burstcount_1(\hps_f2h_sdram0_data_burstcount[1]~input_o ),
	.hps_f2h_sdram0_data_burstcount_2(\hps_f2h_sdram0_data_burstcount[2]~input_o ),
	.hps_f2h_sdram0_data_burstcount_3(\hps_f2h_sdram0_data_burstcount[3]~input_o ),
	.hps_f2h_sdram0_data_burstcount_4(\hps_f2h_sdram0_data_burstcount[4]~input_o ),
	.hps_f2h_sdram0_data_burstcount_5(\hps_f2h_sdram0_data_burstcount[5]~input_o ),
	.hps_f2h_sdram0_data_burstcount_6(\hps_f2h_sdram0_data_burstcount[6]~input_o ),
	.hps_f2h_sdram0_data_burstcount_7(\hps_f2h_sdram0_data_burstcount[7]~input_o ),
	.hps_f2h_sdram0_data_writedata_0(\hps_f2h_sdram0_data_writedata[0]~input_o ),
	.hps_f2h_sdram0_data_writedata_1(\hps_f2h_sdram0_data_writedata[1]~input_o ),
	.hps_f2h_sdram0_data_writedata_2(\hps_f2h_sdram0_data_writedata[2]~input_o ),
	.hps_f2h_sdram0_data_writedata_3(\hps_f2h_sdram0_data_writedata[3]~input_o ),
	.hps_f2h_sdram0_data_writedata_4(\hps_f2h_sdram0_data_writedata[4]~input_o ),
	.hps_f2h_sdram0_data_writedata_5(\hps_f2h_sdram0_data_writedata[5]~input_o ),
	.hps_f2h_sdram0_data_writedata_6(\hps_f2h_sdram0_data_writedata[6]~input_o ),
	.hps_f2h_sdram0_data_writedata_7(\hps_f2h_sdram0_data_writedata[7]~input_o ),
	.hps_f2h_sdram0_data_writedata_8(\hps_f2h_sdram0_data_writedata[8]~input_o ),
	.hps_f2h_sdram0_data_writedata_9(\hps_f2h_sdram0_data_writedata[9]~input_o ),
	.hps_f2h_sdram0_data_writedata_10(\hps_f2h_sdram0_data_writedata[10]~input_o ),
	.hps_f2h_sdram0_data_writedata_11(\hps_f2h_sdram0_data_writedata[11]~input_o ),
	.hps_f2h_sdram0_data_writedata_12(\hps_f2h_sdram0_data_writedata[12]~input_o ),
	.hps_f2h_sdram0_data_writedata_13(\hps_f2h_sdram0_data_writedata[13]~input_o ),
	.hps_f2h_sdram0_data_writedata_14(\hps_f2h_sdram0_data_writedata[14]~input_o ),
	.hps_f2h_sdram0_data_writedata_15(\hps_f2h_sdram0_data_writedata[15]~input_o ),
	.hps_f2h_sdram0_data_writedata_16(\hps_f2h_sdram0_data_writedata[16]~input_o ),
	.hps_f2h_sdram0_data_writedata_17(\hps_f2h_sdram0_data_writedata[17]~input_o ),
	.hps_f2h_sdram0_data_writedata_18(\hps_f2h_sdram0_data_writedata[18]~input_o ),
	.hps_f2h_sdram0_data_writedata_19(\hps_f2h_sdram0_data_writedata[19]~input_o ),
	.hps_f2h_sdram0_data_writedata_20(\hps_f2h_sdram0_data_writedata[20]~input_o ),
	.hps_f2h_sdram0_data_writedata_21(\hps_f2h_sdram0_data_writedata[21]~input_o ),
	.hps_f2h_sdram0_data_writedata_22(\hps_f2h_sdram0_data_writedata[22]~input_o ),
	.hps_f2h_sdram0_data_writedata_23(\hps_f2h_sdram0_data_writedata[23]~input_o ),
	.hps_f2h_sdram0_data_writedata_24(\hps_f2h_sdram0_data_writedata[24]~input_o ),
	.hps_f2h_sdram0_data_writedata_25(\hps_f2h_sdram0_data_writedata[25]~input_o ),
	.hps_f2h_sdram0_data_writedata_26(\hps_f2h_sdram0_data_writedata[26]~input_o ),
	.hps_f2h_sdram0_data_writedata_27(\hps_f2h_sdram0_data_writedata[27]~input_o ),
	.hps_f2h_sdram0_data_writedata_28(\hps_f2h_sdram0_data_writedata[28]~input_o ),
	.hps_f2h_sdram0_data_writedata_29(\hps_f2h_sdram0_data_writedata[29]~input_o ),
	.hps_f2h_sdram0_data_writedata_30(\hps_f2h_sdram0_data_writedata[30]~input_o ),
	.hps_f2h_sdram0_data_writedata_31(\hps_f2h_sdram0_data_writedata[31]~input_o ),
	.hps_f2h_sdram0_data_writedata_32(\hps_f2h_sdram0_data_writedata[32]~input_o ),
	.hps_f2h_sdram0_data_writedata_33(\hps_f2h_sdram0_data_writedata[33]~input_o ),
	.hps_f2h_sdram0_data_writedata_34(\hps_f2h_sdram0_data_writedata[34]~input_o ),
	.hps_f2h_sdram0_data_writedata_35(\hps_f2h_sdram0_data_writedata[35]~input_o ),
	.hps_f2h_sdram0_data_writedata_36(\hps_f2h_sdram0_data_writedata[36]~input_o ),
	.hps_f2h_sdram0_data_writedata_37(\hps_f2h_sdram0_data_writedata[37]~input_o ),
	.hps_f2h_sdram0_data_writedata_38(\hps_f2h_sdram0_data_writedata[38]~input_o ),
	.hps_f2h_sdram0_data_writedata_39(\hps_f2h_sdram0_data_writedata[39]~input_o ),
	.hps_f2h_sdram0_data_writedata_40(\hps_f2h_sdram0_data_writedata[40]~input_o ),
	.hps_f2h_sdram0_data_writedata_41(\hps_f2h_sdram0_data_writedata[41]~input_o ),
	.hps_f2h_sdram0_data_writedata_42(\hps_f2h_sdram0_data_writedata[42]~input_o ),
	.hps_f2h_sdram0_data_writedata_43(\hps_f2h_sdram0_data_writedata[43]~input_o ),
	.hps_f2h_sdram0_data_writedata_44(\hps_f2h_sdram0_data_writedata[44]~input_o ),
	.hps_f2h_sdram0_data_writedata_45(\hps_f2h_sdram0_data_writedata[45]~input_o ),
	.hps_f2h_sdram0_data_writedata_46(\hps_f2h_sdram0_data_writedata[46]~input_o ),
	.hps_f2h_sdram0_data_writedata_47(\hps_f2h_sdram0_data_writedata[47]~input_o ),
	.hps_f2h_sdram0_data_writedata_48(\hps_f2h_sdram0_data_writedata[48]~input_o ),
	.hps_f2h_sdram0_data_writedata_49(\hps_f2h_sdram0_data_writedata[49]~input_o ),
	.hps_f2h_sdram0_data_writedata_50(\hps_f2h_sdram0_data_writedata[50]~input_o ),
	.hps_f2h_sdram0_data_writedata_51(\hps_f2h_sdram0_data_writedata[51]~input_o ),
	.hps_f2h_sdram0_data_writedata_52(\hps_f2h_sdram0_data_writedata[52]~input_o ),
	.hps_f2h_sdram0_data_writedata_53(\hps_f2h_sdram0_data_writedata[53]~input_o ),
	.hps_f2h_sdram0_data_writedata_54(\hps_f2h_sdram0_data_writedata[54]~input_o ),
	.hps_f2h_sdram0_data_writedata_55(\hps_f2h_sdram0_data_writedata[55]~input_o ),
	.hps_f2h_sdram0_data_writedata_56(\hps_f2h_sdram0_data_writedata[56]~input_o ),
	.hps_f2h_sdram0_data_writedata_57(\hps_f2h_sdram0_data_writedata[57]~input_o ),
	.hps_f2h_sdram0_data_writedata_58(\hps_f2h_sdram0_data_writedata[58]~input_o ),
	.hps_f2h_sdram0_data_writedata_59(\hps_f2h_sdram0_data_writedata[59]~input_o ),
	.hps_f2h_sdram0_data_writedata_60(\hps_f2h_sdram0_data_writedata[60]~input_o ),
	.hps_f2h_sdram0_data_writedata_61(\hps_f2h_sdram0_data_writedata[61]~input_o ),
	.hps_f2h_sdram0_data_writedata_62(\hps_f2h_sdram0_data_writedata[62]~input_o ),
	.hps_f2h_sdram0_data_writedata_63(\hps_f2h_sdram0_data_writedata[63]~input_o ),
	.hps_f2h_sdram0_data_byteenable_0(\hps_f2h_sdram0_data_byteenable[0]~input_o ),
	.hps_f2h_sdram0_data_byteenable_1(\hps_f2h_sdram0_data_byteenable[1]~input_o ),
	.hps_f2h_sdram0_data_byteenable_2(\hps_f2h_sdram0_data_byteenable[2]~input_o ),
	.hps_f2h_sdram0_data_byteenable_3(\hps_f2h_sdram0_data_byteenable[3]~input_o ),
	.hps_f2h_sdram0_data_byteenable_4(\hps_f2h_sdram0_data_byteenable[4]~input_o ),
	.hps_f2h_sdram0_data_byteenable_5(\hps_f2h_sdram0_data_byteenable[5]~input_o ),
	.hps_f2h_sdram0_data_byteenable_6(\hps_f2h_sdram0_data_byteenable[6]~input_o ),
	.hps_f2h_sdram0_data_byteenable_7(\hps_f2h_sdram0_data_byteenable[7]~input_o ),
	.hps_f2h_sdram0_data_writedata_64(\hps_f2h_sdram0_data_writedata[64]~input_o ),
	.hps_f2h_sdram0_data_writedata_65(\hps_f2h_sdram0_data_writedata[65]~input_o ),
	.hps_f2h_sdram0_data_writedata_66(\hps_f2h_sdram0_data_writedata[66]~input_o ),
	.hps_f2h_sdram0_data_writedata_67(\hps_f2h_sdram0_data_writedata[67]~input_o ),
	.hps_f2h_sdram0_data_writedata_68(\hps_f2h_sdram0_data_writedata[68]~input_o ),
	.hps_f2h_sdram0_data_writedata_69(\hps_f2h_sdram0_data_writedata[69]~input_o ),
	.hps_f2h_sdram0_data_writedata_70(\hps_f2h_sdram0_data_writedata[70]~input_o ),
	.hps_f2h_sdram0_data_writedata_71(\hps_f2h_sdram0_data_writedata[71]~input_o ),
	.hps_f2h_sdram0_data_writedata_72(\hps_f2h_sdram0_data_writedata[72]~input_o ),
	.hps_f2h_sdram0_data_writedata_73(\hps_f2h_sdram0_data_writedata[73]~input_o ),
	.hps_f2h_sdram0_data_writedata_74(\hps_f2h_sdram0_data_writedata[74]~input_o ),
	.hps_f2h_sdram0_data_writedata_75(\hps_f2h_sdram0_data_writedata[75]~input_o ),
	.hps_f2h_sdram0_data_writedata_76(\hps_f2h_sdram0_data_writedata[76]~input_o ),
	.hps_f2h_sdram0_data_writedata_77(\hps_f2h_sdram0_data_writedata[77]~input_o ),
	.hps_f2h_sdram0_data_writedata_78(\hps_f2h_sdram0_data_writedata[78]~input_o ),
	.hps_f2h_sdram0_data_writedata_79(\hps_f2h_sdram0_data_writedata[79]~input_o ),
	.hps_f2h_sdram0_data_writedata_80(\hps_f2h_sdram0_data_writedata[80]~input_o ),
	.hps_f2h_sdram0_data_writedata_81(\hps_f2h_sdram0_data_writedata[81]~input_o ),
	.hps_f2h_sdram0_data_writedata_82(\hps_f2h_sdram0_data_writedata[82]~input_o ),
	.hps_f2h_sdram0_data_writedata_83(\hps_f2h_sdram0_data_writedata[83]~input_o ),
	.hps_f2h_sdram0_data_writedata_84(\hps_f2h_sdram0_data_writedata[84]~input_o ),
	.hps_f2h_sdram0_data_writedata_85(\hps_f2h_sdram0_data_writedata[85]~input_o ),
	.hps_f2h_sdram0_data_writedata_86(\hps_f2h_sdram0_data_writedata[86]~input_o ),
	.hps_f2h_sdram0_data_writedata_87(\hps_f2h_sdram0_data_writedata[87]~input_o ),
	.hps_f2h_sdram0_data_writedata_88(\hps_f2h_sdram0_data_writedata[88]~input_o ),
	.hps_f2h_sdram0_data_writedata_89(\hps_f2h_sdram0_data_writedata[89]~input_o ),
	.hps_f2h_sdram0_data_writedata_90(\hps_f2h_sdram0_data_writedata[90]~input_o ),
	.hps_f2h_sdram0_data_writedata_91(\hps_f2h_sdram0_data_writedata[91]~input_o ),
	.hps_f2h_sdram0_data_writedata_92(\hps_f2h_sdram0_data_writedata[92]~input_o ),
	.hps_f2h_sdram0_data_writedata_93(\hps_f2h_sdram0_data_writedata[93]~input_o ),
	.hps_f2h_sdram0_data_writedata_94(\hps_f2h_sdram0_data_writedata[94]~input_o ),
	.hps_f2h_sdram0_data_writedata_95(\hps_f2h_sdram0_data_writedata[95]~input_o ),
	.hps_f2h_sdram0_data_writedata_96(\hps_f2h_sdram0_data_writedata[96]~input_o ),
	.hps_f2h_sdram0_data_writedata_97(\hps_f2h_sdram0_data_writedata[97]~input_o ),
	.hps_f2h_sdram0_data_writedata_98(\hps_f2h_sdram0_data_writedata[98]~input_o ),
	.hps_f2h_sdram0_data_writedata_99(\hps_f2h_sdram0_data_writedata[99]~input_o ),
	.hps_f2h_sdram0_data_writedata_100(\hps_f2h_sdram0_data_writedata[100]~input_o ),
	.hps_f2h_sdram0_data_writedata_101(\hps_f2h_sdram0_data_writedata[101]~input_o ),
	.hps_f2h_sdram0_data_writedata_102(\hps_f2h_sdram0_data_writedata[102]~input_o ),
	.hps_f2h_sdram0_data_writedata_103(\hps_f2h_sdram0_data_writedata[103]~input_o ),
	.hps_f2h_sdram0_data_writedata_104(\hps_f2h_sdram0_data_writedata[104]~input_o ),
	.hps_f2h_sdram0_data_writedata_105(\hps_f2h_sdram0_data_writedata[105]~input_o ),
	.hps_f2h_sdram0_data_writedata_106(\hps_f2h_sdram0_data_writedata[106]~input_o ),
	.hps_f2h_sdram0_data_writedata_107(\hps_f2h_sdram0_data_writedata[107]~input_o ),
	.hps_f2h_sdram0_data_writedata_108(\hps_f2h_sdram0_data_writedata[108]~input_o ),
	.hps_f2h_sdram0_data_writedata_109(\hps_f2h_sdram0_data_writedata[109]~input_o ),
	.hps_f2h_sdram0_data_writedata_110(\hps_f2h_sdram0_data_writedata[110]~input_o ),
	.hps_f2h_sdram0_data_writedata_111(\hps_f2h_sdram0_data_writedata[111]~input_o ),
	.hps_f2h_sdram0_data_writedata_112(\hps_f2h_sdram0_data_writedata[112]~input_o ),
	.hps_f2h_sdram0_data_writedata_113(\hps_f2h_sdram0_data_writedata[113]~input_o ),
	.hps_f2h_sdram0_data_writedata_114(\hps_f2h_sdram0_data_writedata[114]~input_o ),
	.hps_f2h_sdram0_data_writedata_115(\hps_f2h_sdram0_data_writedata[115]~input_o ),
	.hps_f2h_sdram0_data_writedata_116(\hps_f2h_sdram0_data_writedata[116]~input_o ),
	.hps_f2h_sdram0_data_writedata_117(\hps_f2h_sdram0_data_writedata[117]~input_o ),
	.hps_f2h_sdram0_data_writedata_118(\hps_f2h_sdram0_data_writedata[118]~input_o ),
	.hps_f2h_sdram0_data_writedata_119(\hps_f2h_sdram0_data_writedata[119]~input_o ),
	.hps_f2h_sdram0_data_writedata_120(\hps_f2h_sdram0_data_writedata[120]~input_o ),
	.hps_f2h_sdram0_data_writedata_121(\hps_f2h_sdram0_data_writedata[121]~input_o ),
	.hps_f2h_sdram0_data_writedata_122(\hps_f2h_sdram0_data_writedata[122]~input_o ),
	.hps_f2h_sdram0_data_writedata_123(\hps_f2h_sdram0_data_writedata[123]~input_o ),
	.hps_f2h_sdram0_data_writedata_124(\hps_f2h_sdram0_data_writedata[124]~input_o ),
	.hps_f2h_sdram0_data_writedata_125(\hps_f2h_sdram0_data_writedata[125]~input_o ),
	.hps_f2h_sdram0_data_writedata_126(\hps_f2h_sdram0_data_writedata[126]~input_o ),
	.hps_f2h_sdram0_data_writedata_127(\hps_f2h_sdram0_data_writedata[127]~input_o ),
	.hps_f2h_sdram0_data_byteenable_8(\hps_f2h_sdram0_data_byteenable[8]~input_o ),
	.hps_f2h_sdram0_data_byteenable_9(\hps_f2h_sdram0_data_byteenable[9]~input_o ),
	.hps_f2h_sdram0_data_byteenable_10(\hps_f2h_sdram0_data_byteenable[10]~input_o ),
	.hps_f2h_sdram0_data_byteenable_11(\hps_f2h_sdram0_data_byteenable[11]~input_o ),
	.hps_f2h_sdram0_data_byteenable_12(\hps_f2h_sdram0_data_byteenable[12]~input_o ),
	.hps_f2h_sdram0_data_byteenable_13(\hps_f2h_sdram0_data_byteenable[13]~input_o ),
	.hps_f2h_sdram0_data_byteenable_14(\hps_f2h_sdram0_data_byteenable[14]~input_o ),
	.hps_f2h_sdram0_data_byteenable_15(\hps_f2h_sdram0_data_byteenable[15]~input_o ),
	.hps_f2h_sdram0_data_writedata_128(\hps_f2h_sdram0_data_writedata[128]~input_o ),
	.hps_f2h_sdram0_data_writedata_129(\hps_f2h_sdram0_data_writedata[129]~input_o ),
	.hps_f2h_sdram0_data_writedata_130(\hps_f2h_sdram0_data_writedata[130]~input_o ),
	.hps_f2h_sdram0_data_writedata_131(\hps_f2h_sdram0_data_writedata[131]~input_o ),
	.hps_f2h_sdram0_data_writedata_132(\hps_f2h_sdram0_data_writedata[132]~input_o ),
	.hps_f2h_sdram0_data_writedata_133(\hps_f2h_sdram0_data_writedata[133]~input_o ),
	.hps_f2h_sdram0_data_writedata_134(\hps_f2h_sdram0_data_writedata[134]~input_o ),
	.hps_f2h_sdram0_data_writedata_135(\hps_f2h_sdram0_data_writedata[135]~input_o ),
	.hps_f2h_sdram0_data_writedata_136(\hps_f2h_sdram0_data_writedata[136]~input_o ),
	.hps_f2h_sdram0_data_writedata_137(\hps_f2h_sdram0_data_writedata[137]~input_o ),
	.hps_f2h_sdram0_data_writedata_138(\hps_f2h_sdram0_data_writedata[138]~input_o ),
	.hps_f2h_sdram0_data_writedata_139(\hps_f2h_sdram0_data_writedata[139]~input_o ),
	.hps_f2h_sdram0_data_writedata_140(\hps_f2h_sdram0_data_writedata[140]~input_o ),
	.hps_f2h_sdram0_data_writedata_141(\hps_f2h_sdram0_data_writedata[141]~input_o ),
	.hps_f2h_sdram0_data_writedata_142(\hps_f2h_sdram0_data_writedata[142]~input_o ),
	.hps_f2h_sdram0_data_writedata_143(\hps_f2h_sdram0_data_writedata[143]~input_o ),
	.hps_f2h_sdram0_data_writedata_144(\hps_f2h_sdram0_data_writedata[144]~input_o ),
	.hps_f2h_sdram0_data_writedata_145(\hps_f2h_sdram0_data_writedata[145]~input_o ),
	.hps_f2h_sdram0_data_writedata_146(\hps_f2h_sdram0_data_writedata[146]~input_o ),
	.hps_f2h_sdram0_data_writedata_147(\hps_f2h_sdram0_data_writedata[147]~input_o ),
	.hps_f2h_sdram0_data_writedata_148(\hps_f2h_sdram0_data_writedata[148]~input_o ),
	.hps_f2h_sdram0_data_writedata_149(\hps_f2h_sdram0_data_writedata[149]~input_o ),
	.hps_f2h_sdram0_data_writedata_150(\hps_f2h_sdram0_data_writedata[150]~input_o ),
	.hps_f2h_sdram0_data_writedata_151(\hps_f2h_sdram0_data_writedata[151]~input_o ),
	.hps_f2h_sdram0_data_writedata_152(\hps_f2h_sdram0_data_writedata[152]~input_o ),
	.hps_f2h_sdram0_data_writedata_153(\hps_f2h_sdram0_data_writedata[153]~input_o ),
	.hps_f2h_sdram0_data_writedata_154(\hps_f2h_sdram0_data_writedata[154]~input_o ),
	.hps_f2h_sdram0_data_writedata_155(\hps_f2h_sdram0_data_writedata[155]~input_o ),
	.hps_f2h_sdram0_data_writedata_156(\hps_f2h_sdram0_data_writedata[156]~input_o ),
	.hps_f2h_sdram0_data_writedata_157(\hps_f2h_sdram0_data_writedata[157]~input_o ),
	.hps_f2h_sdram0_data_writedata_158(\hps_f2h_sdram0_data_writedata[158]~input_o ),
	.hps_f2h_sdram0_data_writedata_159(\hps_f2h_sdram0_data_writedata[159]~input_o ),
	.hps_f2h_sdram0_data_writedata_160(\hps_f2h_sdram0_data_writedata[160]~input_o ),
	.hps_f2h_sdram0_data_writedata_161(\hps_f2h_sdram0_data_writedata[161]~input_o ),
	.hps_f2h_sdram0_data_writedata_162(\hps_f2h_sdram0_data_writedata[162]~input_o ),
	.hps_f2h_sdram0_data_writedata_163(\hps_f2h_sdram0_data_writedata[163]~input_o ),
	.hps_f2h_sdram0_data_writedata_164(\hps_f2h_sdram0_data_writedata[164]~input_o ),
	.hps_f2h_sdram0_data_writedata_165(\hps_f2h_sdram0_data_writedata[165]~input_o ),
	.hps_f2h_sdram0_data_writedata_166(\hps_f2h_sdram0_data_writedata[166]~input_o ),
	.hps_f2h_sdram0_data_writedata_167(\hps_f2h_sdram0_data_writedata[167]~input_o ),
	.hps_f2h_sdram0_data_writedata_168(\hps_f2h_sdram0_data_writedata[168]~input_o ),
	.hps_f2h_sdram0_data_writedata_169(\hps_f2h_sdram0_data_writedata[169]~input_o ),
	.hps_f2h_sdram0_data_writedata_170(\hps_f2h_sdram0_data_writedata[170]~input_o ),
	.hps_f2h_sdram0_data_writedata_171(\hps_f2h_sdram0_data_writedata[171]~input_o ),
	.hps_f2h_sdram0_data_writedata_172(\hps_f2h_sdram0_data_writedata[172]~input_o ),
	.hps_f2h_sdram0_data_writedata_173(\hps_f2h_sdram0_data_writedata[173]~input_o ),
	.hps_f2h_sdram0_data_writedata_174(\hps_f2h_sdram0_data_writedata[174]~input_o ),
	.hps_f2h_sdram0_data_writedata_175(\hps_f2h_sdram0_data_writedata[175]~input_o ),
	.hps_f2h_sdram0_data_writedata_176(\hps_f2h_sdram0_data_writedata[176]~input_o ),
	.hps_f2h_sdram0_data_writedata_177(\hps_f2h_sdram0_data_writedata[177]~input_o ),
	.hps_f2h_sdram0_data_writedata_178(\hps_f2h_sdram0_data_writedata[178]~input_o ),
	.hps_f2h_sdram0_data_writedata_179(\hps_f2h_sdram0_data_writedata[179]~input_o ),
	.hps_f2h_sdram0_data_writedata_180(\hps_f2h_sdram0_data_writedata[180]~input_o ),
	.hps_f2h_sdram0_data_writedata_181(\hps_f2h_sdram0_data_writedata[181]~input_o ),
	.hps_f2h_sdram0_data_writedata_182(\hps_f2h_sdram0_data_writedata[182]~input_o ),
	.hps_f2h_sdram0_data_writedata_183(\hps_f2h_sdram0_data_writedata[183]~input_o ),
	.hps_f2h_sdram0_data_writedata_184(\hps_f2h_sdram0_data_writedata[184]~input_o ),
	.hps_f2h_sdram0_data_writedata_185(\hps_f2h_sdram0_data_writedata[185]~input_o ),
	.hps_f2h_sdram0_data_writedata_186(\hps_f2h_sdram0_data_writedata[186]~input_o ),
	.hps_f2h_sdram0_data_writedata_187(\hps_f2h_sdram0_data_writedata[187]~input_o ),
	.hps_f2h_sdram0_data_writedata_188(\hps_f2h_sdram0_data_writedata[188]~input_o ),
	.hps_f2h_sdram0_data_writedata_189(\hps_f2h_sdram0_data_writedata[189]~input_o ),
	.hps_f2h_sdram0_data_writedata_190(\hps_f2h_sdram0_data_writedata[190]~input_o ),
	.hps_f2h_sdram0_data_writedata_191(\hps_f2h_sdram0_data_writedata[191]~input_o ),
	.hps_f2h_sdram0_data_byteenable_16(\hps_f2h_sdram0_data_byteenable[16]~input_o ),
	.hps_f2h_sdram0_data_byteenable_17(\hps_f2h_sdram0_data_byteenable[17]~input_o ),
	.hps_f2h_sdram0_data_byteenable_18(\hps_f2h_sdram0_data_byteenable[18]~input_o ),
	.hps_f2h_sdram0_data_byteenable_19(\hps_f2h_sdram0_data_byteenable[19]~input_o ),
	.hps_f2h_sdram0_data_byteenable_20(\hps_f2h_sdram0_data_byteenable[20]~input_o ),
	.hps_f2h_sdram0_data_byteenable_21(\hps_f2h_sdram0_data_byteenable[21]~input_o ),
	.hps_f2h_sdram0_data_byteenable_22(\hps_f2h_sdram0_data_byteenable[22]~input_o ),
	.hps_f2h_sdram0_data_byteenable_23(\hps_f2h_sdram0_data_byteenable[23]~input_o ),
	.hps_f2h_sdram0_data_writedata_192(\hps_f2h_sdram0_data_writedata[192]~input_o ),
	.hps_f2h_sdram0_data_writedata_193(\hps_f2h_sdram0_data_writedata[193]~input_o ),
	.hps_f2h_sdram0_data_writedata_194(\hps_f2h_sdram0_data_writedata[194]~input_o ),
	.hps_f2h_sdram0_data_writedata_195(\hps_f2h_sdram0_data_writedata[195]~input_o ),
	.hps_f2h_sdram0_data_writedata_196(\hps_f2h_sdram0_data_writedata[196]~input_o ),
	.hps_f2h_sdram0_data_writedata_197(\hps_f2h_sdram0_data_writedata[197]~input_o ),
	.hps_f2h_sdram0_data_writedata_198(\hps_f2h_sdram0_data_writedata[198]~input_o ),
	.hps_f2h_sdram0_data_writedata_199(\hps_f2h_sdram0_data_writedata[199]~input_o ),
	.hps_f2h_sdram0_data_writedata_200(\hps_f2h_sdram0_data_writedata[200]~input_o ),
	.hps_f2h_sdram0_data_writedata_201(\hps_f2h_sdram0_data_writedata[201]~input_o ),
	.hps_f2h_sdram0_data_writedata_202(\hps_f2h_sdram0_data_writedata[202]~input_o ),
	.hps_f2h_sdram0_data_writedata_203(\hps_f2h_sdram0_data_writedata[203]~input_o ),
	.hps_f2h_sdram0_data_writedata_204(\hps_f2h_sdram0_data_writedata[204]~input_o ),
	.hps_f2h_sdram0_data_writedata_205(\hps_f2h_sdram0_data_writedata[205]~input_o ),
	.hps_f2h_sdram0_data_writedata_206(\hps_f2h_sdram0_data_writedata[206]~input_o ),
	.hps_f2h_sdram0_data_writedata_207(\hps_f2h_sdram0_data_writedata[207]~input_o ),
	.hps_f2h_sdram0_data_writedata_208(\hps_f2h_sdram0_data_writedata[208]~input_o ),
	.hps_f2h_sdram0_data_writedata_209(\hps_f2h_sdram0_data_writedata[209]~input_o ),
	.hps_f2h_sdram0_data_writedata_210(\hps_f2h_sdram0_data_writedata[210]~input_o ),
	.hps_f2h_sdram0_data_writedata_211(\hps_f2h_sdram0_data_writedata[211]~input_o ),
	.hps_f2h_sdram0_data_writedata_212(\hps_f2h_sdram0_data_writedata[212]~input_o ),
	.hps_f2h_sdram0_data_writedata_213(\hps_f2h_sdram0_data_writedata[213]~input_o ),
	.hps_f2h_sdram0_data_writedata_214(\hps_f2h_sdram0_data_writedata[214]~input_o ),
	.hps_f2h_sdram0_data_writedata_215(\hps_f2h_sdram0_data_writedata[215]~input_o ),
	.hps_f2h_sdram0_data_writedata_216(\hps_f2h_sdram0_data_writedata[216]~input_o ),
	.hps_f2h_sdram0_data_writedata_217(\hps_f2h_sdram0_data_writedata[217]~input_o ),
	.hps_f2h_sdram0_data_writedata_218(\hps_f2h_sdram0_data_writedata[218]~input_o ),
	.hps_f2h_sdram0_data_writedata_219(\hps_f2h_sdram0_data_writedata[219]~input_o ),
	.hps_f2h_sdram0_data_writedata_220(\hps_f2h_sdram0_data_writedata[220]~input_o ),
	.hps_f2h_sdram0_data_writedata_221(\hps_f2h_sdram0_data_writedata[221]~input_o ),
	.hps_f2h_sdram0_data_writedata_222(\hps_f2h_sdram0_data_writedata[222]~input_o ),
	.hps_f2h_sdram0_data_writedata_223(\hps_f2h_sdram0_data_writedata[223]~input_o ),
	.hps_f2h_sdram0_data_writedata_224(\hps_f2h_sdram0_data_writedata[224]~input_o ),
	.hps_f2h_sdram0_data_writedata_225(\hps_f2h_sdram0_data_writedata[225]~input_o ),
	.hps_f2h_sdram0_data_writedata_226(\hps_f2h_sdram0_data_writedata[226]~input_o ),
	.hps_f2h_sdram0_data_writedata_227(\hps_f2h_sdram0_data_writedata[227]~input_o ),
	.hps_f2h_sdram0_data_writedata_228(\hps_f2h_sdram0_data_writedata[228]~input_o ),
	.hps_f2h_sdram0_data_writedata_229(\hps_f2h_sdram0_data_writedata[229]~input_o ),
	.hps_f2h_sdram0_data_writedata_230(\hps_f2h_sdram0_data_writedata[230]~input_o ),
	.hps_f2h_sdram0_data_writedata_231(\hps_f2h_sdram0_data_writedata[231]~input_o ),
	.hps_f2h_sdram0_data_writedata_232(\hps_f2h_sdram0_data_writedata[232]~input_o ),
	.hps_f2h_sdram0_data_writedata_233(\hps_f2h_sdram0_data_writedata[233]~input_o ),
	.hps_f2h_sdram0_data_writedata_234(\hps_f2h_sdram0_data_writedata[234]~input_o ),
	.hps_f2h_sdram0_data_writedata_235(\hps_f2h_sdram0_data_writedata[235]~input_o ),
	.hps_f2h_sdram0_data_writedata_236(\hps_f2h_sdram0_data_writedata[236]~input_o ),
	.hps_f2h_sdram0_data_writedata_237(\hps_f2h_sdram0_data_writedata[237]~input_o ),
	.hps_f2h_sdram0_data_writedata_238(\hps_f2h_sdram0_data_writedata[238]~input_o ),
	.hps_f2h_sdram0_data_writedata_239(\hps_f2h_sdram0_data_writedata[239]~input_o ),
	.hps_f2h_sdram0_data_writedata_240(\hps_f2h_sdram0_data_writedata[240]~input_o ),
	.hps_f2h_sdram0_data_writedata_241(\hps_f2h_sdram0_data_writedata[241]~input_o ),
	.hps_f2h_sdram0_data_writedata_242(\hps_f2h_sdram0_data_writedata[242]~input_o ),
	.hps_f2h_sdram0_data_writedata_243(\hps_f2h_sdram0_data_writedata[243]~input_o ),
	.hps_f2h_sdram0_data_writedata_244(\hps_f2h_sdram0_data_writedata[244]~input_o ),
	.hps_f2h_sdram0_data_writedata_245(\hps_f2h_sdram0_data_writedata[245]~input_o ),
	.hps_f2h_sdram0_data_writedata_246(\hps_f2h_sdram0_data_writedata[246]~input_o ),
	.hps_f2h_sdram0_data_writedata_247(\hps_f2h_sdram0_data_writedata[247]~input_o ),
	.hps_f2h_sdram0_data_writedata_248(\hps_f2h_sdram0_data_writedata[248]~input_o ),
	.hps_f2h_sdram0_data_writedata_249(\hps_f2h_sdram0_data_writedata[249]~input_o ),
	.hps_f2h_sdram0_data_writedata_250(\hps_f2h_sdram0_data_writedata[250]~input_o ),
	.hps_f2h_sdram0_data_writedata_251(\hps_f2h_sdram0_data_writedata[251]~input_o ),
	.hps_f2h_sdram0_data_writedata_252(\hps_f2h_sdram0_data_writedata[252]~input_o ),
	.hps_f2h_sdram0_data_writedata_253(\hps_f2h_sdram0_data_writedata[253]~input_o ),
	.hps_f2h_sdram0_data_writedata_254(\hps_f2h_sdram0_data_writedata[254]~input_o ),
	.hps_f2h_sdram0_data_writedata_255(\hps_f2h_sdram0_data_writedata[255]~input_o ),
	.hps_f2h_sdram0_data_byteenable_24(\hps_f2h_sdram0_data_byteenable[24]~input_o ),
	.hps_f2h_sdram0_data_byteenable_25(\hps_f2h_sdram0_data_byteenable[25]~input_o ),
	.hps_f2h_sdram0_data_byteenable_26(\hps_f2h_sdram0_data_byteenable[26]~input_o ),
	.hps_f2h_sdram0_data_byteenable_27(\hps_f2h_sdram0_data_byteenable[27]~input_o ),
	.hps_f2h_sdram0_data_byteenable_28(\hps_f2h_sdram0_data_byteenable[28]~input_o ),
	.hps_f2h_sdram0_data_byteenable_29(\hps_f2h_sdram0_data_byteenable[29]~input_o ),
	.hps_f2h_sdram0_data_byteenable_30(\hps_f2h_sdram0_data_byteenable[30]~input_o ),
	.hps_f2h_sdram0_data_byteenable_31(\hps_f2h_sdram0_data_byteenable[31]~input_o ));

terminal_qsys_terminal_qsys_base_address_ddr_1 control(
	.data_out_0(\control|data_out[0]~q ),
	.data_out_1(\control|data_out[1]~q ),
	.data_out_2(\control|data_out[2]~q ),
	.data_out_3(\control|data_out[3]~q ),
	.data_out_4(\control|data_out[4]~q ),
	.data_out_5(\control|data_out[5]~q ),
	.data_out_6(\control|data_out[6]~q ),
	.data_out_7(\control|data_out[7]~q ),
	.data_out_8(\control|data_out[8]~q ),
	.data_out_9(\control|data_out[9]~q ),
	.data_out_10(\control|data_out[10]~q ),
	.data_out_11(\control|data_out[11]~q ),
	.data_out_12(\control|data_out[12]~q ),
	.data_out_13(\control|data_out[13]~q ),
	.data_out_14(\control|data_out[14]~q ),
	.data_out_15(\control|data_out[15]~q ),
	.data_out_16(\control|data_out[16]~q ),
	.data_out_17(\control|data_out[17]~q ),
	.data_out_18(\control|data_out[18]~q ),
	.data_out_19(\control|data_out[19]~q ),
	.data_out_20(\control|data_out[20]~q ),
	.data_out_21(\control|data_out[21]~q ),
	.data_out_22(\control|data_out[22]~q ),
	.data_out_23(\control|data_out[23]~q ),
	.data_out_24(\control|data_out[24]~q ),
	.data_out_25(\control|data_out[25]~q ),
	.data_out_26(\control|data_out[26]~q ),
	.data_out_27(\control|data_out[27]~q ),
	.data_out_28(\control|data_out[28]~q ),
	.data_out_29(\control|data_out[29]~q ),
	.data_out_30(\control|data_out[30]~q ),
	.data_out_31(\control|data_out[31]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|control_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|control_s1_translator|wait_latency_counter[0]~q ),
	.writedata({\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ,
\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ,\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q }),
	.reset_n(\rst_controller_001|rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|control_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\control|readdata[0]~combout ),
	.readdata_1(\control|readdata[1]~combout ),
	.readdata_2(\control|readdata[2]~combout ),
	.readdata_3(\control|readdata[3]~combout ),
	.readdata_4(\control|readdata[4]~combout ),
	.readdata_5(\control|readdata[5]~combout ),
	.readdata_6(\control|readdata[6]~combout ),
	.readdata_7(\control|readdata[7]~combout ),
	.readdata_8(\control|readdata[8]~combout ),
	.readdata_9(\control|readdata[9]~combout ),
	.readdata_10(\control|readdata[10]~combout ),
	.readdata_11(\control|readdata[11]~combout ),
	.readdata_12(\control|readdata[12]~combout ),
	.readdata_13(\control|readdata[13]~combout ),
	.readdata_14(\control|readdata[14]~combout ),
	.readdata_15(\control|readdata[15]~combout ),
	.readdata_16(\control|readdata[16]~combout ),
	.readdata_17(\control|readdata[17]~combout ),
	.readdata_18(\control|readdata[18]~combout ),
	.readdata_19(\control|readdata[19]~combout ),
	.readdata_20(\control|readdata[20]~combout ),
	.readdata_21(\control|readdata[21]~combout ),
	.readdata_22(\control|readdata[22]~combout ),
	.readdata_23(\control|readdata[23]~combout ),
	.readdata_24(\control|readdata[24]~combout ),
	.readdata_25(\control|readdata[25]~combout ),
	.readdata_26(\control|readdata[26]~combout ),
	.readdata_27(\control|readdata[27]~combout ),
	.readdata_28(\control|readdata[28]~combout ),
	.readdata_29(\control|readdata[29]~combout ),
	.readdata_30(\control|readdata[30]~combout ),
	.readdata_31(\control|readdata[31]~combout ),
	.clk(\clk_clk~input_o ));

terminal_qsys_terminal_qsys_base_address_ddr base_address_ddr(
	.data_out_0(\base_address_ddr|data_out[0]~q ),
	.data_out_1(\base_address_ddr|data_out[1]~q ),
	.data_out_2(\base_address_ddr|data_out[2]~q ),
	.data_out_3(\base_address_ddr|data_out[3]~q ),
	.data_out_4(\base_address_ddr|data_out[4]~q ),
	.data_out_5(\base_address_ddr|data_out[5]~q ),
	.data_out_6(\base_address_ddr|data_out[6]~q ),
	.data_out_7(\base_address_ddr|data_out[7]~q ),
	.data_out_8(\base_address_ddr|data_out[8]~q ),
	.data_out_9(\base_address_ddr|data_out[9]~q ),
	.data_out_10(\base_address_ddr|data_out[10]~q ),
	.data_out_11(\base_address_ddr|data_out[11]~q ),
	.data_out_12(\base_address_ddr|data_out[12]~q ),
	.data_out_13(\base_address_ddr|data_out[13]~q ),
	.data_out_14(\base_address_ddr|data_out[14]~q ),
	.data_out_15(\base_address_ddr|data_out[15]~q ),
	.data_out_16(\base_address_ddr|data_out[16]~q ),
	.data_out_17(\base_address_ddr|data_out[17]~q ),
	.data_out_18(\base_address_ddr|data_out[18]~q ),
	.data_out_19(\base_address_ddr|data_out[19]~q ),
	.data_out_20(\base_address_ddr|data_out[20]~q ),
	.data_out_21(\base_address_ddr|data_out[21]~q ),
	.data_out_22(\base_address_ddr|data_out[22]~q ),
	.data_out_23(\base_address_ddr|data_out[23]~q ),
	.data_out_24(\base_address_ddr|data_out[24]~q ),
	.data_out_25(\base_address_ddr|data_out[25]~q ),
	.data_out_26(\base_address_ddr|data_out[26]~q ),
	.data_out_27(\base_address_ddr|data_out[27]~q ),
	.data_out_28(\base_address_ddr|data_out[28]~q ),
	.data_out_29(\base_address_ddr|data_out[29]~q ),
	.data_out_30(\base_address_ddr|data_out[30]~q ),
	.data_out_31(\base_address_ddr|data_out[31]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|base_address_ddr_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|base_address_ddr_s1_translator|wait_latency_counter[0]~q ),
	.writedata({\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ,
\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ,\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q }),
	.reset_n(\rst_controller|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|base_address_ddr_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\base_address_ddr|readdata[0]~combout ),
	.readdata_1(\base_address_ddr|readdata[1]~combout ),
	.readdata_2(\base_address_ddr|readdata[2]~combout ),
	.readdata_3(\base_address_ddr|readdata[3]~combout ),
	.readdata_4(\base_address_ddr|readdata[4]~combout ),
	.readdata_5(\base_address_ddr|readdata[5]~combout ),
	.readdata_6(\base_address_ddr|readdata[6]~combout ),
	.readdata_7(\base_address_ddr|readdata[7]~combout ),
	.readdata_8(\base_address_ddr|readdata[8]~combout ),
	.readdata_9(\base_address_ddr|readdata[9]~combout ),
	.readdata_10(\base_address_ddr|readdata[10]~combout ),
	.readdata_11(\base_address_ddr|readdata[11]~combout ),
	.readdata_12(\base_address_ddr|readdata[12]~combout ),
	.readdata_13(\base_address_ddr|readdata[13]~combout ),
	.readdata_14(\base_address_ddr|readdata[14]~combout ),
	.readdata_15(\base_address_ddr|readdata[15]~combout ),
	.readdata_16(\base_address_ddr|readdata[16]~combout ),
	.readdata_17(\base_address_ddr|readdata[17]~combout ),
	.readdata_18(\base_address_ddr|readdata[18]~combout ),
	.readdata_19(\base_address_ddr|readdata[19]~combout ),
	.readdata_20(\base_address_ddr|readdata[20]~combout ),
	.readdata_21(\base_address_ddr|readdata[21]~combout ),
	.readdata_22(\base_address_ddr|readdata[22]~combout ),
	.readdata_23(\base_address_ddr|readdata[23]~combout ),
	.readdata_24(\base_address_ddr|readdata[24]~combout ),
	.readdata_25(\base_address_ddr|readdata[25]~combout ),
	.readdata_26(\base_address_ddr|readdata[26]~combout ),
	.readdata_27(\base_address_ddr|readdata[27]~combout ),
	.readdata_28(\base_address_ddr|readdata[28]~combout ),
	.readdata_29(\base_address_ddr|readdata[29]~combout ),
	.readdata_30(\base_address_ddr|readdata[30]~combout ),
	.readdata_31(\base_address_ddr|readdata[31]~combout ),
	.clk(\clk_clk~input_o ));

terminal_qsys_terminal_qsys_mm_interconnect_0 mm_interconnect_0(
	.h2f_lw_ARVALID_0(\hps|fpga_interfaces|h2f_lw_ARVALID[0] ),
	.h2f_lw_AWVALID_0(\hps|fpga_interfaces|h2f_lw_AWVALID[0] ),
	.h2f_lw_BREADY_0(\hps|fpga_interfaces|h2f_lw_BREADY[0] ),
	.h2f_lw_RREADY_0(\hps|fpga_interfaces|h2f_lw_RREADY[0] ),
	.h2f_lw_WLAST_0(\hps|fpga_interfaces|h2f_lw_WLAST[0] ),
	.h2f_lw_WVALID_0(\hps|fpga_interfaces|h2f_lw_WVALID[0] ),
	.h2f_lw_ARADDR_0(\hps|fpga_interfaces|h2f_lw_ARADDR[0] ),
	.h2f_lw_ARADDR_1(\hps|fpga_interfaces|h2f_lw_ARADDR[1] ),
	.h2f_lw_ARADDR_2(\hps|fpga_interfaces|h2f_lw_ARADDR[2] ),
	.h2f_lw_ARADDR_3(\hps|fpga_interfaces|h2f_lw_ARADDR[3] ),
	.h2f_lw_ARADDR_4(\hps|fpga_interfaces|h2f_lw_ARADDR[4] ),
	.h2f_lw_ARADDR_5(\hps|fpga_interfaces|h2f_lw_ARADDR[5] ),
	.h2f_lw_ARADDR_6(\hps|fpga_interfaces|h2f_lw_ARADDR[6] ),
	.h2f_lw_ARADDR_7(\hps|fpga_interfaces|h2f_lw_ARADDR[7] ),
	.h2f_lw_ARADDR_8(\hps|fpga_interfaces|h2f_lw_ARADDR[8] ),
	.h2f_lw_ARADDR_9(\hps|fpga_interfaces|h2f_lw_ARADDR[9] ),
	.h2f_lw_ARADDR_10(\hps|fpga_interfaces|h2f_lw_ARADDR[10] ),
	.h2f_lw_ARADDR_11(\hps|fpga_interfaces|h2f_lw_ARADDR[11] ),
	.h2f_lw_ARADDR_12(\hps|fpga_interfaces|h2f_lw_ARADDR[12] ),
	.h2f_lw_ARADDR_13(\hps|fpga_interfaces|h2f_lw_ARADDR[13] ),
	.h2f_lw_ARADDR_14(\hps|fpga_interfaces|h2f_lw_ARADDR[14] ),
	.h2f_lw_ARADDR_15(\hps|fpga_interfaces|h2f_lw_ARADDR[15] ),
	.h2f_lw_ARADDR_16(\hps|fpga_interfaces|h2f_lw_ARADDR[16] ),
	.h2f_lw_ARADDR_17(\hps|fpga_interfaces|h2f_lw_ARADDR[17] ),
	.h2f_lw_ARADDR_18(\hps|fpga_interfaces|h2f_lw_ARADDR[18] ),
	.h2f_lw_ARBURST_0(\hps|fpga_interfaces|h2f_lw_ARBURST[0] ),
	.h2f_lw_ARBURST_1(\hps|fpga_interfaces|h2f_lw_ARBURST[1] ),
	.h2f_lw_ARID_0(\hps|fpga_interfaces|h2f_lw_ARID[0] ),
	.h2f_lw_ARID_1(\hps|fpga_interfaces|h2f_lw_ARID[1] ),
	.h2f_lw_ARID_2(\hps|fpga_interfaces|h2f_lw_ARID[2] ),
	.h2f_lw_ARID_3(\hps|fpga_interfaces|h2f_lw_ARID[3] ),
	.h2f_lw_ARID_4(\hps|fpga_interfaces|h2f_lw_ARID[4] ),
	.h2f_lw_ARID_5(\hps|fpga_interfaces|h2f_lw_ARID[5] ),
	.h2f_lw_ARID_6(\hps|fpga_interfaces|h2f_lw_ARID[6] ),
	.h2f_lw_ARID_7(\hps|fpga_interfaces|h2f_lw_ARID[7] ),
	.h2f_lw_ARID_8(\hps|fpga_interfaces|h2f_lw_ARID[8] ),
	.h2f_lw_ARID_9(\hps|fpga_interfaces|h2f_lw_ARID[9] ),
	.h2f_lw_ARID_10(\hps|fpga_interfaces|h2f_lw_ARID[10] ),
	.h2f_lw_ARID_11(\hps|fpga_interfaces|h2f_lw_ARID[11] ),
	.h2f_lw_ARLEN_0(\hps|fpga_interfaces|h2f_lw_ARLEN[0] ),
	.h2f_lw_ARLEN_1(\hps|fpga_interfaces|h2f_lw_ARLEN[1] ),
	.h2f_lw_ARLEN_2(\hps|fpga_interfaces|h2f_lw_ARLEN[2] ),
	.h2f_lw_ARLEN_3(\hps|fpga_interfaces|h2f_lw_ARLEN[3] ),
	.h2f_lw_ARSIZE_0(\hps|fpga_interfaces|h2f_lw_ARSIZE[0] ),
	.h2f_lw_ARSIZE_1(\hps|fpga_interfaces|h2f_lw_ARSIZE[1] ),
	.h2f_lw_ARSIZE_2(\hps|fpga_interfaces|h2f_lw_ARSIZE[2] ),
	.h2f_lw_AWADDR_0(\hps|fpga_interfaces|h2f_lw_AWADDR[0] ),
	.h2f_lw_AWADDR_1(\hps|fpga_interfaces|h2f_lw_AWADDR[1] ),
	.h2f_lw_AWADDR_2(\hps|fpga_interfaces|h2f_lw_AWADDR[2] ),
	.h2f_lw_AWADDR_3(\hps|fpga_interfaces|h2f_lw_AWADDR[3] ),
	.h2f_lw_AWADDR_4(\hps|fpga_interfaces|h2f_lw_AWADDR[4] ),
	.h2f_lw_AWADDR_5(\hps|fpga_interfaces|h2f_lw_AWADDR[5] ),
	.h2f_lw_AWADDR_6(\hps|fpga_interfaces|h2f_lw_AWADDR[6] ),
	.h2f_lw_AWADDR_7(\hps|fpga_interfaces|h2f_lw_AWADDR[7] ),
	.h2f_lw_AWADDR_8(\hps|fpga_interfaces|h2f_lw_AWADDR[8] ),
	.h2f_lw_AWADDR_9(\hps|fpga_interfaces|h2f_lw_AWADDR[9] ),
	.h2f_lw_AWADDR_10(\hps|fpga_interfaces|h2f_lw_AWADDR[10] ),
	.h2f_lw_AWADDR_11(\hps|fpga_interfaces|h2f_lw_AWADDR[11] ),
	.h2f_lw_AWADDR_12(\hps|fpga_interfaces|h2f_lw_AWADDR[12] ),
	.h2f_lw_AWADDR_13(\hps|fpga_interfaces|h2f_lw_AWADDR[13] ),
	.h2f_lw_AWADDR_14(\hps|fpga_interfaces|h2f_lw_AWADDR[14] ),
	.h2f_lw_AWADDR_15(\hps|fpga_interfaces|h2f_lw_AWADDR[15] ),
	.h2f_lw_AWADDR_16(\hps|fpga_interfaces|h2f_lw_AWADDR[16] ),
	.h2f_lw_AWADDR_17(\hps|fpga_interfaces|h2f_lw_AWADDR[17] ),
	.h2f_lw_AWADDR_18(\hps|fpga_interfaces|h2f_lw_AWADDR[18] ),
	.h2f_lw_AWBURST_0(\hps|fpga_interfaces|h2f_lw_AWBURST[0] ),
	.h2f_lw_AWBURST_1(\hps|fpga_interfaces|h2f_lw_AWBURST[1] ),
	.h2f_lw_AWID_0(\hps|fpga_interfaces|h2f_lw_AWID[0] ),
	.h2f_lw_AWID_1(\hps|fpga_interfaces|h2f_lw_AWID[1] ),
	.h2f_lw_AWID_2(\hps|fpga_interfaces|h2f_lw_AWID[2] ),
	.h2f_lw_AWID_3(\hps|fpga_interfaces|h2f_lw_AWID[3] ),
	.h2f_lw_AWID_4(\hps|fpga_interfaces|h2f_lw_AWID[4] ),
	.h2f_lw_AWID_5(\hps|fpga_interfaces|h2f_lw_AWID[5] ),
	.h2f_lw_AWID_6(\hps|fpga_interfaces|h2f_lw_AWID[6] ),
	.h2f_lw_AWID_7(\hps|fpga_interfaces|h2f_lw_AWID[7] ),
	.h2f_lw_AWID_8(\hps|fpga_interfaces|h2f_lw_AWID[8] ),
	.h2f_lw_AWID_9(\hps|fpga_interfaces|h2f_lw_AWID[9] ),
	.h2f_lw_AWID_10(\hps|fpga_interfaces|h2f_lw_AWID[10] ),
	.h2f_lw_AWID_11(\hps|fpga_interfaces|h2f_lw_AWID[11] ),
	.h2f_lw_AWLEN_0(\hps|fpga_interfaces|h2f_lw_AWLEN[0] ),
	.h2f_lw_AWLEN_1(\hps|fpga_interfaces|h2f_lw_AWLEN[1] ),
	.h2f_lw_AWLEN_2(\hps|fpga_interfaces|h2f_lw_AWLEN[2] ),
	.h2f_lw_AWLEN_3(\hps|fpga_interfaces|h2f_lw_AWLEN[3] ),
	.h2f_lw_AWSIZE_0(\hps|fpga_interfaces|h2f_lw_AWSIZE[0] ),
	.h2f_lw_AWSIZE_1(\hps|fpga_interfaces|h2f_lw_AWSIZE[1] ),
	.h2f_lw_AWSIZE_2(\hps|fpga_interfaces|h2f_lw_AWSIZE[2] ),
	.h2f_lw_WDATA_0(\hps|fpga_interfaces|h2f_lw_WDATA[0] ),
	.h2f_lw_WDATA_1(\hps|fpga_interfaces|h2f_lw_WDATA[1] ),
	.h2f_lw_WDATA_2(\hps|fpga_interfaces|h2f_lw_WDATA[2] ),
	.h2f_lw_WDATA_3(\hps|fpga_interfaces|h2f_lw_WDATA[3] ),
	.h2f_lw_WDATA_4(\hps|fpga_interfaces|h2f_lw_WDATA[4] ),
	.h2f_lw_WDATA_5(\hps|fpga_interfaces|h2f_lw_WDATA[5] ),
	.h2f_lw_WDATA_6(\hps|fpga_interfaces|h2f_lw_WDATA[6] ),
	.h2f_lw_WDATA_7(\hps|fpga_interfaces|h2f_lw_WDATA[7] ),
	.h2f_lw_WDATA_8(\hps|fpga_interfaces|h2f_lw_WDATA[8] ),
	.h2f_lw_WDATA_9(\hps|fpga_interfaces|h2f_lw_WDATA[9] ),
	.h2f_lw_WDATA_10(\hps|fpga_interfaces|h2f_lw_WDATA[10] ),
	.h2f_lw_WDATA_11(\hps|fpga_interfaces|h2f_lw_WDATA[11] ),
	.h2f_lw_WDATA_12(\hps|fpga_interfaces|h2f_lw_WDATA[12] ),
	.h2f_lw_WDATA_13(\hps|fpga_interfaces|h2f_lw_WDATA[13] ),
	.h2f_lw_WDATA_14(\hps|fpga_interfaces|h2f_lw_WDATA[14] ),
	.h2f_lw_WDATA_15(\hps|fpga_interfaces|h2f_lw_WDATA[15] ),
	.h2f_lw_WDATA_16(\hps|fpga_interfaces|h2f_lw_WDATA[16] ),
	.h2f_lw_WDATA_17(\hps|fpga_interfaces|h2f_lw_WDATA[17] ),
	.h2f_lw_WDATA_18(\hps|fpga_interfaces|h2f_lw_WDATA[18] ),
	.h2f_lw_WDATA_19(\hps|fpga_interfaces|h2f_lw_WDATA[19] ),
	.h2f_lw_WDATA_20(\hps|fpga_interfaces|h2f_lw_WDATA[20] ),
	.h2f_lw_WDATA_21(\hps|fpga_interfaces|h2f_lw_WDATA[21] ),
	.h2f_lw_WDATA_22(\hps|fpga_interfaces|h2f_lw_WDATA[22] ),
	.h2f_lw_WDATA_23(\hps|fpga_interfaces|h2f_lw_WDATA[23] ),
	.h2f_lw_WDATA_24(\hps|fpga_interfaces|h2f_lw_WDATA[24] ),
	.h2f_lw_WDATA_25(\hps|fpga_interfaces|h2f_lw_WDATA[25] ),
	.h2f_lw_WDATA_26(\hps|fpga_interfaces|h2f_lw_WDATA[26] ),
	.h2f_lw_WDATA_27(\hps|fpga_interfaces|h2f_lw_WDATA[27] ),
	.h2f_lw_WDATA_28(\hps|fpga_interfaces|h2f_lw_WDATA[28] ),
	.h2f_lw_WDATA_29(\hps|fpga_interfaces|h2f_lw_WDATA[29] ),
	.h2f_lw_WDATA_30(\hps|fpga_interfaces|h2f_lw_WDATA[30] ),
	.h2f_lw_WDATA_31(\hps|fpga_interfaces|h2f_lw_WDATA[31] ),
	.h2f_lw_WSTRB_0(\hps|fpga_interfaces|h2f_lw_WSTRB[0] ),
	.h2f_lw_WSTRB_1(\hps|fpga_interfaces|h2f_lw_WSTRB[1] ),
	.h2f_lw_WSTRB_2(\hps|fpga_interfaces|h2f_lw_WSTRB[2] ),
	.h2f_lw_WSTRB_3(\hps|fpga_interfaces|h2f_lw_WSTRB[3] ),
	.wait_latency_counter_1(\mm_interconnect_0|base_address_ddr_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|base_address_ddr_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_11(\mm_interconnect_0|control_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|control_s1_translator|wait_latency_counter[0]~q ),
	.wait_latency_counter_12(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_02(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[0]~q ),
	.cmd_sink_ready(\mm_interconnect_0|hps_h2f_lw_axi_master_rd_limiter|cmd_sink_ready~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload_0(\mm_interconnect_0|rsp_mux_001|src_payload[0]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.nonposted_cmd_accepted1(\mm_interconnect_0|hps_h2f_lw_axi_master_wr_limiter|nonposted_cmd_accepted~1_combout ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux_001|src_data[0]~5_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux_001|src_data[1]~11_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux_001|src_data[2]~17_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux_001|src_data[3]~23_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux_001|src_data[4]~29_combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux_001|src_data[5]~35_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux_001|src_data[6]~41_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux_001|src_data[7]~48_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux_001|src_data[8]~54_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux_001|src_data[9]~58_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux_001|src_payload~11_combout ),
	.src_payload13(\mm_interconnect_0|rsp_mux_001|src_payload~14_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux_001|src_payload~17_combout ),
	.src_payload15(\mm_interconnect_0|rsp_mux_001|src_payload~20_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux_001|src_payload~23_combout ),
	.src_payload17(\mm_interconnect_0|rsp_mux_001|src_payload~26_combout ),
	.src_payload18(\mm_interconnect_0|rsp_mux_001|src_payload~29_combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux_001|src_payload~32_combout ),
	.src_payload20(\mm_interconnect_0|rsp_mux_001|src_payload~35_combout ),
	.src_payload21(\mm_interconnect_0|rsp_mux_001|src_payload~38_combout ),
	.src_payload22(\mm_interconnect_0|rsp_mux_001|src_payload~41_combout ),
	.src_payload23(\mm_interconnect_0|rsp_mux_001|src_payload~44_combout ),
	.src_payload24(\mm_interconnect_0|rsp_mux_001|src_payload~47_combout ),
	.src_payload25(\mm_interconnect_0|rsp_mux_001|src_payload~50_combout ),
	.src_payload26(\mm_interconnect_0|rsp_mux_001|src_payload~53_combout ),
	.src_payload27(\mm_interconnect_0|rsp_mux_001|src_payload~56_combout ),
	.src_payload28(\mm_interconnect_0|rsp_mux_001|src_payload~59_combout ),
	.src_payload29(\mm_interconnect_0|rsp_mux_001|src_payload~62_combout ),
	.src_payload30(\mm_interconnect_0|rsp_mux_001|src_payload~65_combout ),
	.src_payload31(\mm_interconnect_0|rsp_mux_001|src_payload~68_combout ),
	.src_payload32(\mm_interconnect_0|rsp_mux_001|src_payload~71_combout ),
	.src_payload33(\mm_interconnect_0|rsp_mux_001|src_payload~74_combout ),
	.src_data_92(\mm_interconnect_0|rsp_mux_001|src_data[92]~combout ),
	.src_data_93(\mm_interconnect_0|rsp_mux_001|src_data[93]~combout ),
	.src_data_94(\mm_interconnect_0|rsp_mux_001|src_data[94]~combout ),
	.src_data_95(\mm_interconnect_0|rsp_mux_001|src_data[95]~combout ),
	.src_data_96(\mm_interconnect_0|rsp_mux_001|src_data[96]~combout ),
	.src_data_97(\mm_interconnect_0|rsp_mux_001|src_data[97]~combout ),
	.src_data_98(\mm_interconnect_0|rsp_mux_001|src_data[98]~combout ),
	.src_data_99(\mm_interconnect_0|rsp_mux_001|src_data[99]~combout ),
	.src_data_100(\mm_interconnect_0|rsp_mux_001|src_data[100]~combout ),
	.src_data_101(\mm_interconnect_0|rsp_mux_001|src_data[101]~combout ),
	.src_data_102(\mm_interconnect_0|rsp_mux_001|src_data[102]~combout ),
	.src_data_103(\mm_interconnect_0|rsp_mux_001|src_data[103]~combout ),
	.in_data_reg_0(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write(\mm_interconnect_0|base_address_ddr_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_1(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_2(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_3(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_4(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_5(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_6(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_7(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_8(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_9(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_10(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_11(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_12(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_13(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_14(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_15(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_16(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_17(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_18(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_19(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_20(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_21(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_22(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_23(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_24(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_25(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_26(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_27(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_28(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_29(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_30(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_31(\mm_interconnect_0|base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.in_data_reg_01(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.altera_reset_synchronizer_int_chain_out1(\rst_controller_001|rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.m0_write1(\mm_interconnect_0|control_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_31(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_21(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_110(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_210(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_32(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_41(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_51(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_61(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_71(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_81(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_91(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.in_data_reg_101(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[10]~q ),
	.in_data_reg_111(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[11]~q ),
	.in_data_reg_121(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[12]~q ),
	.in_data_reg_131(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[13]~q ),
	.in_data_reg_141(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[14]~q ),
	.in_data_reg_151(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[15]~q ),
	.in_data_reg_161(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[16]~q ),
	.in_data_reg_171(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[17]~q ),
	.in_data_reg_181(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[18]~q ),
	.in_data_reg_191(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[19]~q ),
	.in_data_reg_201(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[20]~q ),
	.in_data_reg_211(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[21]~q ),
	.in_data_reg_221(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[22]~q ),
	.in_data_reg_231(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[23]~q ),
	.in_data_reg_241(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[24]~q ),
	.in_data_reg_251(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[25]~q ),
	.in_data_reg_261(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[26]~q ),
	.in_data_reg_271(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[27]~q ),
	.in_data_reg_281(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[28]~q ),
	.in_data_reg_291(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[29]~q ),
	.in_data_reg_301(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[30]~q ),
	.in_data_reg_311(\mm_interconnect_0|control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[31]~q ),
	.in_data_reg_02(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q ),
	.m0_write2(\mm_interconnect_0|leds_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_32(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_22(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_112(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ),
	.in_data_reg_212(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ),
	.in_data_reg_33(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ),
	.in_data_reg_42(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ),
	.in_data_reg_52(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ),
	.in_data_reg_62(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ),
	.in_data_reg_72(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ),
	.in_data_reg_82(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ),
	.in_data_reg_92(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ),
	.altera_reset_synchronizer_int_chain_out2(\rst_controller_002|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\control|readdata[0]~combout ),
	.readdata_01(\base_address_ddr|readdata[0]~combout ),
	.readdata_02(\leds|readdata[0]~combout ),
	.readdata_03(\state|readdata[0]~q ),
	.readdata_04(\switches|readdata[0]~q ),
	.readdata_1(\control|readdata[1]~combout ),
	.readdata_11(\base_address_ddr|readdata[1]~combout ),
	.readdata_12(\leds|readdata[1]~combout ),
	.readdata_13(\state|readdata[1]~q ),
	.readdata_14(\switches|readdata[1]~q ),
	.readdata_2(\control|readdata[2]~combout ),
	.readdata_21(\base_address_ddr|readdata[2]~combout ),
	.readdata_22(\leds|readdata[2]~combout ),
	.readdata_23(\state|readdata[2]~q ),
	.readdata_24(\switches|readdata[2]~q ),
	.readdata_3(\control|readdata[3]~combout ),
	.readdata_31(\base_address_ddr|readdata[3]~combout ),
	.readdata_32(\leds|readdata[3]~combout ),
	.readdata_33(\state|readdata[3]~q ),
	.readdata_34(\switches|readdata[3]~q ),
	.readdata_4(\control|readdata[4]~combout ),
	.readdata_41(\base_address_ddr|readdata[4]~combout ),
	.readdata_42(\leds|readdata[4]~combout ),
	.readdata_43(\state|readdata[4]~q ),
	.readdata_44(\switches|readdata[4]~q ),
	.readdata_5(\control|readdata[5]~combout ),
	.readdata_51(\base_address_ddr|readdata[5]~combout ),
	.readdata_52(\leds|readdata[5]~combout ),
	.readdata_53(\state|readdata[5]~q ),
	.readdata_54(\switches|readdata[5]~q ),
	.readdata_6(\control|readdata[6]~combout ),
	.readdata_61(\base_address_ddr|readdata[6]~combout ),
	.readdata_62(\leds|readdata[6]~combout ),
	.readdata_63(\state|readdata[6]~q ),
	.readdata_64(\switches|readdata[6]~q ),
	.readdata_7(\control|readdata[7]~combout ),
	.readdata_71(\base_address_ddr|readdata[7]~combout ),
	.readdata_72(\leds|readdata[7]~combout ),
	.readdata_73(\state|readdata[7]~q ),
	.readdata_74(\switches|readdata[7]~q ),
	.readdata_8(\control|readdata[8]~combout ),
	.readdata_81(\base_address_ddr|readdata[8]~combout ),
	.readdata_82(\leds|readdata[8]~combout ),
	.readdata_83(\state|readdata[8]~q ),
	.readdata_84(\switches|readdata[8]~q ),
	.readdata_9(\state|readdata[9]~q ),
	.readdata_91(\control|readdata[9]~combout ),
	.readdata_92(\base_address_ddr|readdata[9]~combout ),
	.readdata_93(\leds|readdata[9]~combout ),
	.readdata_94(\switches|readdata[9]~q ),
	.readdata_10(\control|readdata[10]~combout ),
	.readdata_101(\base_address_ddr|readdata[10]~combout ),
	.readdata_102(\state|readdata[10]~q ),
	.readdata_111(\control|readdata[11]~combout ),
	.readdata_112(\base_address_ddr|readdata[11]~combout ),
	.readdata_113(\state|readdata[11]~q ),
	.readdata_121(\base_address_ddr|readdata[12]~combout ),
	.readdata_122(\control|readdata[12]~combout ),
	.readdata_123(\state|readdata[12]~q ),
	.readdata_131(\base_address_ddr|readdata[13]~combout ),
	.readdata_132(\control|readdata[13]~combout ),
	.readdata_133(\state|readdata[13]~q ),
	.readdata_141(\base_address_ddr|readdata[14]~combout ),
	.readdata_142(\control|readdata[14]~combout ),
	.readdata_143(\state|readdata[14]~q ),
	.readdata_15(\base_address_ddr|readdata[15]~combout ),
	.readdata_151(\control|readdata[15]~combout ),
	.readdata_152(\state|readdata[15]~q ),
	.readdata_16(\base_address_ddr|readdata[16]~combout ),
	.readdata_161(\control|readdata[16]~combout ),
	.readdata_162(\state|readdata[16]~q ),
	.readdata_17(\base_address_ddr|readdata[17]~combout ),
	.readdata_171(\control|readdata[17]~combout ),
	.readdata_172(\state|readdata[17]~q ),
	.readdata_18(\base_address_ddr|readdata[18]~combout ),
	.readdata_181(\control|readdata[18]~combout ),
	.readdata_182(\state|readdata[18]~q ),
	.readdata_19(\control|readdata[19]~combout ),
	.readdata_191(\base_address_ddr|readdata[19]~combout ),
	.readdata_192(\state|readdata[19]~q ),
	.readdata_20(\control|readdata[20]~combout ),
	.readdata_201(\base_address_ddr|readdata[20]~combout ),
	.readdata_202(\state|readdata[20]~q ),
	.readdata_211(\control|readdata[21]~combout ),
	.readdata_212(\base_address_ddr|readdata[21]~combout ),
	.readdata_213(\state|readdata[21]~q ),
	.readdata_221(\base_address_ddr|readdata[22]~combout ),
	.readdata_222(\control|readdata[22]~combout ),
	.readdata_223(\state|readdata[22]~q ),
	.readdata_231(\base_address_ddr|readdata[23]~combout ),
	.readdata_232(\control|readdata[23]~combout ),
	.readdata_233(\state|readdata[23]~q ),
	.readdata_241(\control|readdata[24]~combout ),
	.readdata_242(\base_address_ddr|readdata[24]~combout ),
	.readdata_243(\state|readdata[24]~q ),
	.readdata_25(\base_address_ddr|readdata[25]~combout ),
	.readdata_251(\control|readdata[25]~combout ),
	.readdata_252(\state|readdata[25]~q ),
	.readdata_26(\base_address_ddr|readdata[26]~combout ),
	.readdata_261(\control|readdata[26]~combout ),
	.readdata_262(\state|readdata[26]~q ),
	.readdata_27(\control|readdata[27]~combout ),
	.readdata_271(\base_address_ddr|readdata[27]~combout ),
	.readdata_272(\state|readdata[27]~q ),
	.readdata_28(\control|readdata[28]~combout ),
	.readdata_281(\base_address_ddr|readdata[28]~combout ),
	.readdata_282(\state|readdata[28]~q ),
	.readdata_29(\base_address_ddr|readdata[29]~combout ),
	.readdata_291(\control|readdata[29]~combout ),
	.readdata_292(\state|readdata[29]~q ),
	.readdata_30(\control|readdata[30]~combout ),
	.readdata_301(\base_address_ddr|readdata[30]~combout ),
	.readdata_302(\state|readdata[30]~q ),
	.readdata_311(\base_address_ddr|readdata[31]~combout ),
	.readdata_312(\control|readdata[31]~combout ),
	.readdata_313(\state|readdata[31]~q ),
	.int_nxt_addr_reg_dly_33(\mm_interconnect_0|state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_23(\mm_interconnect_0|state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.int_nxt_addr_reg_dly_34(\mm_interconnect_0|switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_24(\mm_interconnect_0|switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ));

terminal_qsys_terminal_qsys_switches switches(
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\switches|readdata[0]~q ),
	.readdata_1(\switches|readdata[1]~q ),
	.readdata_2(\switches|readdata[2]~q ),
	.readdata_3(\switches|readdata[3]~q ),
	.readdata_4(\switches|readdata[4]~q ),
	.readdata_5(\switches|readdata[5]~q ),
	.readdata_6(\switches|readdata[6]~q ),
	.readdata_7(\switches|readdata[7]~q ),
	.readdata_8(\switches|readdata[8]~q ),
	.readdata_9(\switches|readdata[9]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.switches_in_export_0(\switches_in_export[0]~input_o ),
	.switches_in_export_1(\switches_in_export[1]~input_o ),
	.switches_in_export_2(\switches_in_export[2]~input_o ),
	.switches_in_export_3(\switches_in_export[3]~input_o ),
	.switches_in_export_4(\switches_in_export[4]~input_o ),
	.switches_in_export_5(\switches_in_export[5]~input_o ),
	.switches_in_export_6(\switches_in_export[6]~input_o ),
	.switches_in_export_7(\switches_in_export[7]~input_o ),
	.switches_in_export_8(\switches_in_export[8]~input_o ),
	.switches_in_export_9(\switches_in_export[9]~input_o ));

terminal_qsys_terminal_qsys_state state(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.readdata_0(\state|readdata[0]~q ),
	.readdata_1(\state|readdata[1]~q ),
	.readdata_2(\state|readdata[2]~q ),
	.readdata_3(\state|readdata[3]~q ),
	.readdata_4(\state|readdata[4]~q ),
	.readdata_5(\state|readdata[5]~q ),
	.readdata_6(\state|readdata[6]~q ),
	.readdata_7(\state|readdata[7]~q ),
	.readdata_8(\state|readdata[8]~q ),
	.readdata_9(\state|readdata[9]~q ),
	.readdata_10(\state|readdata[10]~q ),
	.readdata_11(\state|readdata[11]~q ),
	.readdata_12(\state|readdata[12]~q ),
	.readdata_13(\state|readdata[13]~q ),
	.readdata_14(\state|readdata[14]~q ),
	.readdata_15(\state|readdata[15]~q ),
	.readdata_16(\state|readdata[16]~q ),
	.readdata_17(\state|readdata[17]~q ),
	.readdata_18(\state|readdata[18]~q ),
	.readdata_19(\state|readdata[19]~q ),
	.readdata_20(\state|readdata[20]~q ),
	.readdata_21(\state|readdata[21]~q ),
	.readdata_22(\state|readdata[22]~q ),
	.readdata_23(\state|readdata[23]~q ),
	.readdata_24(\state|readdata[24]~q ),
	.readdata_25(\state|readdata[25]~q ),
	.readdata_26(\state|readdata[26]~q ),
	.readdata_27(\state|readdata[27]~q ),
	.readdata_28(\state|readdata[28]~q ),
	.readdata_29(\state|readdata[29]~q ),
	.readdata_30(\state|readdata[30]~q ),
	.readdata_31(\state|readdata[31]~q ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.state_in_export_0(\state_in_export[0]~input_o ),
	.state_in_export_1(\state_in_export[1]~input_o ),
	.state_in_export_2(\state_in_export[2]~input_o ),
	.state_in_export_3(\state_in_export[3]~input_o ),
	.state_in_export_4(\state_in_export[4]~input_o ),
	.state_in_export_5(\state_in_export[5]~input_o ),
	.state_in_export_6(\state_in_export[6]~input_o ),
	.state_in_export_7(\state_in_export[7]~input_o ),
	.state_in_export_8(\state_in_export[8]~input_o ),
	.state_in_export_9(\state_in_export[9]~input_o ),
	.state_in_export_10(\state_in_export[10]~input_o ),
	.state_in_export_11(\state_in_export[11]~input_o ),
	.state_in_export_12(\state_in_export[12]~input_o ),
	.state_in_export_13(\state_in_export[13]~input_o ),
	.state_in_export_14(\state_in_export[14]~input_o ),
	.state_in_export_15(\state_in_export[15]~input_o ),
	.state_in_export_16(\state_in_export[16]~input_o ),
	.state_in_export_17(\state_in_export[17]~input_o ),
	.state_in_export_18(\state_in_export[18]~input_o ),
	.state_in_export_19(\state_in_export[19]~input_o ),
	.state_in_export_20(\state_in_export[20]~input_o ),
	.state_in_export_21(\state_in_export[21]~input_o ),
	.state_in_export_22(\state_in_export[22]~input_o ),
	.state_in_export_23(\state_in_export[23]~input_o ),
	.state_in_export_24(\state_in_export[24]~input_o ),
	.state_in_export_25(\state_in_export[25]~input_o ),
	.state_in_export_26(\state_in_export[26]~input_o ),
	.state_in_export_27(\state_in_export[27]~input_o ),
	.state_in_export_28(\state_in_export[28]~input_o ),
	.state_in_export_29(\state_in_export[29]~input_o ),
	.state_in_export_30(\state_in_export[30]~input_o ),
	.state_in_export_31(\state_in_export[31]~input_o ));

terminal_qsys_terminal_qsys_leds leds(
	.data_out_0(\leds|data_out[0]~q ),
	.data_out_1(\leds|data_out[1]~q ),
	.data_out_2(\leds|data_out[2]~q ),
	.data_out_3(\leds|data_out[3]~q ),
	.data_out_4(\leds|data_out[4]~q ),
	.data_out_5(\leds|data_out[5]~q ),
	.data_out_6(\leds|data_out[6]~q ),
	.data_out_7(\leds|data_out[7]~q ),
	.data_out_8(\leds|data_out[8]~q ),
	.data_out_9(\leds|data_out[9]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|leds_s1_translator|wait_latency_counter[0]~q ),
	.reset_n(\rst_controller_001|rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[9]~q ,
\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[8]~q ,\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[7]~q ,
\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[6]~q ,\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[5]~q ,
\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[4]~q ,\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[3]~q ,
\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[2]~q ,\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[1]~q ,
\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[0]~q }),
	.m0_write(\mm_interconnect_0|leds_s1_agent|m0_write~combout ),
	.int_nxt_addr_reg_dly_3(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[3]~q ),
	.int_nxt_addr_reg_dly_2(\mm_interconnect_0|leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.readdata_0(\leds|readdata[0]~combout ),
	.readdata_1(\leds|readdata[1]~combout ),
	.readdata_2(\leds|readdata[2]~combout ),
	.readdata_3(\leds|readdata[3]~combout ),
	.readdata_4(\leds|readdata[4]~combout ),
	.readdata_5(\leds|readdata[5]~combout ),
	.readdata_6(\leds|readdata[6]~combout ),
	.readdata_7(\leds|readdata[7]~combout ),
	.readdata_8(\leds|readdata[8]~combout ),
	.readdata_9(\leds|readdata[9]~combout ),
	.clk(\clk_clk~input_o ));

terminal_qsys_terminal_qsys_rst_controller_1 rst_controller_002(
	.h2f_rst_n_0(\hps|fpga_interfaces|h2f_rst_n[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_002|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ));

terminal_qsys_terminal_qsys_rst_controller_001 rst_controller_001(
	.h2f_rst_n_0(\hps|fpga_interfaces|h2f_rst_n[0] ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller_001|rst_controller_001|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

terminal_qsys_terminal_qsys_rst_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[3]),
	.ibar(memory_mem_dqs_n[3]),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[24]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[25]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[26]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[27]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[28]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[29]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[30]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[31]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[2]),
	.ibar(memory_mem_dqs_n[2]),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[16]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[17]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[18]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[19]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[20]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[21]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[22]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[23]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[1]),
	.ibar(memory_mem_dqs_n[1]),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[8]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[9]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[10]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[11]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[12]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[13]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[14]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[15]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in (
	.i(memory_mem_dqs[0]),
	.ibar(memory_mem_dqs_n[0]),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|dqsin ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .differential_mode = "true";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|strobe_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in (
	.i(memory_mem_dq[0]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in (
	.i(memory_mem_dq[1]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in (
	.i(memory_mem_dq[2]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in (
	.i(memory_mem_dq[3]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in (
	.i(memory_mem_dq[4]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in (
	.i(memory_mem_dq[5]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in (
	.i(memory_mem_dq[6]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_in .simulate_z_as = "z";

cyclonev_io_ibuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in (
	.i(memory_mem_dq[7]),
	.ibar(gnd),
	.dynamicterminationcontrol(gnd),
	.o(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].raw_input ));
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_in .simulate_z_as = "z";

assign \hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~input_o  = hps_hps_io_hps_io_emac1_inst_MDIO;

assign \hps|hps_io|border|hps_io_sdio_inst_CMD[0]~input_o  = hps_hps_io_hps_io_sdio_inst_CMD;

assign \hps|hps_io|border|hps_io_sdio_inst_D0[0]~input_o  = hps_hps_io_hps_io_sdio_inst_D0;

assign \hps|hps_io|border|hps_io_sdio_inst_D1[0]~input_o  = hps_hps_io_hps_io_sdio_inst_D1;

assign \hps|hps_io|border|hps_io_sdio_inst_D2[0]~input_o  = hps_hps_io_hps_io_sdio_inst_D2;

assign \hps|hps_io|border|hps_io_sdio_inst_D3[0]~input_o  = hps_hps_io_hps_io_sdio_inst_D3;

assign \hps_f2h_stm_hw_events_stm_hwevents[0]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[0];

assign \hps_f2h_stm_hw_events_stm_hwevents[1]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[1];

assign \hps_f2h_stm_hw_events_stm_hwevents[2]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[2];

assign \hps_f2h_stm_hw_events_stm_hwevents[3]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[3];

assign \hps_f2h_stm_hw_events_stm_hwevents[4]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[4];

assign \hps_f2h_stm_hw_events_stm_hwevents[5]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[5];

assign \hps_f2h_stm_hw_events_stm_hwevents[6]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[6];

assign \hps_f2h_stm_hw_events_stm_hwevents[7]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[7];

assign \hps_f2h_stm_hw_events_stm_hwevents[8]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[8];

assign \hps_f2h_stm_hw_events_stm_hwevents[9]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[9];

assign \hps_f2h_stm_hw_events_stm_hwevents[10]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[10];

assign \hps_f2h_stm_hw_events_stm_hwevents[11]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[11];

assign \hps_f2h_stm_hw_events_stm_hwevents[12]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[12];

assign \hps_f2h_stm_hw_events_stm_hwevents[13]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[13];

assign \hps_f2h_stm_hw_events_stm_hwevents[14]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[14];

assign \hps_f2h_stm_hw_events_stm_hwevents[15]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[15];

assign \hps_f2h_stm_hw_events_stm_hwevents[16]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[16];

assign \hps_f2h_stm_hw_events_stm_hwevents[17]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[17];

assign \hps_f2h_stm_hw_events_stm_hwevents[18]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[18];

assign \hps_f2h_stm_hw_events_stm_hwevents[19]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[19];

assign \hps_f2h_stm_hw_events_stm_hwevents[20]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[20];

assign \hps_f2h_stm_hw_events_stm_hwevents[21]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[21];

assign \hps_f2h_stm_hw_events_stm_hwevents[22]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[22];

assign \hps_f2h_stm_hw_events_stm_hwevents[23]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[23];

assign \hps_f2h_stm_hw_events_stm_hwevents[24]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[24];

assign \hps_f2h_stm_hw_events_stm_hwevents[25]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[25];

assign \hps_f2h_stm_hw_events_stm_hwevents[26]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[26];

assign \hps_f2h_stm_hw_events_stm_hwevents[27]~input_o  = hps_f2h_stm_hw_events_stm_hwevents[27];

assign \clk_clk~input_o  = clk_clk;

assign \hps_hps_io_hps_io_emac1_inst_RXD0~input_o  = hps_hps_io_hps_io_emac1_inst_RXD0;

assign \hps_hps_io_hps_io_emac1_inst_RXD1~input_o  = hps_hps_io_hps_io_emac1_inst_RXD1;

assign \hps_hps_io_hps_io_emac1_inst_RXD2~input_o  = hps_hps_io_hps_io_emac1_inst_RXD2;

assign \hps_hps_io_hps_io_emac1_inst_RXD3~input_o  = hps_hps_io_hps_io_emac1_inst_RXD3;

assign \hps_hps_io_hps_io_emac1_inst_RX_CLK~input_o  = hps_hps_io_hps_io_emac1_inst_RX_CLK;

assign \hps_hps_io_hps_io_emac1_inst_RX_CTL~input_o  = hps_hps_io_hps_io_emac1_inst_RX_CTL;

assign \hps_hps_io_hps_io_uart0_inst_RX~input_o  = hps_hps_io_hps_io_uart0_inst_RX;

assign \memory_oct_rzqin~input_o  = memory_oct_rzqin;

assign \hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n~input_o  = hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n;

assign \hps_f2h_sdram0_data_read~input_o  = hps_f2h_sdram0_data_read;

assign \hps_f2h_sdram0_data_write~input_o  = hps_f2h_sdram0_data_write;

assign \hps_f2h_sdram0_data_address[0]~input_o  = hps_f2h_sdram0_data_address[0];

assign \hps_f2h_sdram0_data_address[1]~input_o  = hps_f2h_sdram0_data_address[1];

assign \hps_f2h_sdram0_data_address[2]~input_o  = hps_f2h_sdram0_data_address[2];

assign \hps_f2h_sdram0_data_address[3]~input_o  = hps_f2h_sdram0_data_address[3];

assign \hps_f2h_sdram0_data_address[4]~input_o  = hps_f2h_sdram0_data_address[4];

assign \hps_f2h_sdram0_data_address[5]~input_o  = hps_f2h_sdram0_data_address[5];

assign \hps_f2h_sdram0_data_address[6]~input_o  = hps_f2h_sdram0_data_address[6];

assign \hps_f2h_sdram0_data_address[7]~input_o  = hps_f2h_sdram0_data_address[7];

assign \hps_f2h_sdram0_data_address[8]~input_o  = hps_f2h_sdram0_data_address[8];

assign \hps_f2h_sdram0_data_address[9]~input_o  = hps_f2h_sdram0_data_address[9];

assign \hps_f2h_sdram0_data_address[10]~input_o  = hps_f2h_sdram0_data_address[10];

assign \hps_f2h_sdram0_data_address[11]~input_o  = hps_f2h_sdram0_data_address[11];

assign \hps_f2h_sdram0_data_address[12]~input_o  = hps_f2h_sdram0_data_address[12];

assign \hps_f2h_sdram0_data_address[13]~input_o  = hps_f2h_sdram0_data_address[13];

assign \hps_f2h_sdram0_data_address[14]~input_o  = hps_f2h_sdram0_data_address[14];

assign \hps_f2h_sdram0_data_address[15]~input_o  = hps_f2h_sdram0_data_address[15];

assign \hps_f2h_sdram0_data_address[16]~input_o  = hps_f2h_sdram0_data_address[16];

assign \hps_f2h_sdram0_data_address[17]~input_o  = hps_f2h_sdram0_data_address[17];

assign \hps_f2h_sdram0_data_address[18]~input_o  = hps_f2h_sdram0_data_address[18];

assign \hps_f2h_sdram0_data_address[19]~input_o  = hps_f2h_sdram0_data_address[19];

assign \hps_f2h_sdram0_data_address[20]~input_o  = hps_f2h_sdram0_data_address[20];

assign \hps_f2h_sdram0_data_address[21]~input_o  = hps_f2h_sdram0_data_address[21];

assign \hps_f2h_sdram0_data_address[22]~input_o  = hps_f2h_sdram0_data_address[22];

assign \hps_f2h_sdram0_data_address[23]~input_o  = hps_f2h_sdram0_data_address[23];

assign \hps_f2h_sdram0_data_address[24]~input_o  = hps_f2h_sdram0_data_address[24];

assign \hps_f2h_sdram0_data_address[25]~input_o  = hps_f2h_sdram0_data_address[25];

assign \hps_f2h_sdram0_data_address[26]~input_o  = hps_f2h_sdram0_data_address[26];

assign \hps_f2h_sdram0_data_burstcount[0]~input_o  = hps_f2h_sdram0_data_burstcount[0];

assign \hps_f2h_sdram0_data_burstcount[1]~input_o  = hps_f2h_sdram0_data_burstcount[1];

assign \hps_f2h_sdram0_data_burstcount[2]~input_o  = hps_f2h_sdram0_data_burstcount[2];

assign \hps_f2h_sdram0_data_burstcount[3]~input_o  = hps_f2h_sdram0_data_burstcount[3];

assign \hps_f2h_sdram0_data_burstcount[4]~input_o  = hps_f2h_sdram0_data_burstcount[4];

assign \hps_f2h_sdram0_data_burstcount[5]~input_o  = hps_f2h_sdram0_data_burstcount[5];

assign \hps_f2h_sdram0_data_burstcount[6]~input_o  = hps_f2h_sdram0_data_burstcount[6];

assign \hps_f2h_sdram0_data_burstcount[7]~input_o  = hps_f2h_sdram0_data_burstcount[7];

assign \hps_f2h_sdram0_data_writedata[0]~input_o  = hps_f2h_sdram0_data_writedata[0];

assign \hps_f2h_sdram0_data_writedata[1]~input_o  = hps_f2h_sdram0_data_writedata[1];

assign \hps_f2h_sdram0_data_writedata[2]~input_o  = hps_f2h_sdram0_data_writedata[2];

assign \hps_f2h_sdram0_data_writedata[3]~input_o  = hps_f2h_sdram0_data_writedata[3];

assign \hps_f2h_sdram0_data_writedata[4]~input_o  = hps_f2h_sdram0_data_writedata[4];

assign \hps_f2h_sdram0_data_writedata[5]~input_o  = hps_f2h_sdram0_data_writedata[5];

assign \hps_f2h_sdram0_data_writedata[6]~input_o  = hps_f2h_sdram0_data_writedata[6];

assign \hps_f2h_sdram0_data_writedata[7]~input_o  = hps_f2h_sdram0_data_writedata[7];

assign \hps_f2h_sdram0_data_writedata[8]~input_o  = hps_f2h_sdram0_data_writedata[8];

assign \hps_f2h_sdram0_data_writedata[9]~input_o  = hps_f2h_sdram0_data_writedata[9];

assign \hps_f2h_sdram0_data_writedata[10]~input_o  = hps_f2h_sdram0_data_writedata[10];

assign \hps_f2h_sdram0_data_writedata[11]~input_o  = hps_f2h_sdram0_data_writedata[11];

assign \hps_f2h_sdram0_data_writedata[12]~input_o  = hps_f2h_sdram0_data_writedata[12];

assign \hps_f2h_sdram0_data_writedata[13]~input_o  = hps_f2h_sdram0_data_writedata[13];

assign \hps_f2h_sdram0_data_writedata[14]~input_o  = hps_f2h_sdram0_data_writedata[14];

assign \hps_f2h_sdram0_data_writedata[15]~input_o  = hps_f2h_sdram0_data_writedata[15];

assign \hps_f2h_sdram0_data_writedata[16]~input_o  = hps_f2h_sdram0_data_writedata[16];

assign \hps_f2h_sdram0_data_writedata[17]~input_o  = hps_f2h_sdram0_data_writedata[17];

assign \hps_f2h_sdram0_data_writedata[18]~input_o  = hps_f2h_sdram0_data_writedata[18];

assign \hps_f2h_sdram0_data_writedata[19]~input_o  = hps_f2h_sdram0_data_writedata[19];

assign \hps_f2h_sdram0_data_writedata[20]~input_o  = hps_f2h_sdram0_data_writedata[20];

assign \hps_f2h_sdram0_data_writedata[21]~input_o  = hps_f2h_sdram0_data_writedata[21];

assign \hps_f2h_sdram0_data_writedata[22]~input_o  = hps_f2h_sdram0_data_writedata[22];

assign \hps_f2h_sdram0_data_writedata[23]~input_o  = hps_f2h_sdram0_data_writedata[23];

assign \hps_f2h_sdram0_data_writedata[24]~input_o  = hps_f2h_sdram0_data_writedata[24];

assign \hps_f2h_sdram0_data_writedata[25]~input_o  = hps_f2h_sdram0_data_writedata[25];

assign \hps_f2h_sdram0_data_writedata[26]~input_o  = hps_f2h_sdram0_data_writedata[26];

assign \hps_f2h_sdram0_data_writedata[27]~input_o  = hps_f2h_sdram0_data_writedata[27];

assign \hps_f2h_sdram0_data_writedata[28]~input_o  = hps_f2h_sdram0_data_writedata[28];

assign \hps_f2h_sdram0_data_writedata[29]~input_o  = hps_f2h_sdram0_data_writedata[29];

assign \hps_f2h_sdram0_data_writedata[30]~input_o  = hps_f2h_sdram0_data_writedata[30];

assign \hps_f2h_sdram0_data_writedata[31]~input_o  = hps_f2h_sdram0_data_writedata[31];

assign \hps_f2h_sdram0_data_writedata[32]~input_o  = hps_f2h_sdram0_data_writedata[32];

assign \hps_f2h_sdram0_data_writedata[33]~input_o  = hps_f2h_sdram0_data_writedata[33];

assign \hps_f2h_sdram0_data_writedata[34]~input_o  = hps_f2h_sdram0_data_writedata[34];

assign \hps_f2h_sdram0_data_writedata[35]~input_o  = hps_f2h_sdram0_data_writedata[35];

assign \hps_f2h_sdram0_data_writedata[36]~input_o  = hps_f2h_sdram0_data_writedata[36];

assign \hps_f2h_sdram0_data_writedata[37]~input_o  = hps_f2h_sdram0_data_writedata[37];

assign \hps_f2h_sdram0_data_writedata[38]~input_o  = hps_f2h_sdram0_data_writedata[38];

assign \hps_f2h_sdram0_data_writedata[39]~input_o  = hps_f2h_sdram0_data_writedata[39];

assign \hps_f2h_sdram0_data_writedata[40]~input_o  = hps_f2h_sdram0_data_writedata[40];

assign \hps_f2h_sdram0_data_writedata[41]~input_o  = hps_f2h_sdram0_data_writedata[41];

assign \hps_f2h_sdram0_data_writedata[42]~input_o  = hps_f2h_sdram0_data_writedata[42];

assign \hps_f2h_sdram0_data_writedata[43]~input_o  = hps_f2h_sdram0_data_writedata[43];

assign \hps_f2h_sdram0_data_writedata[44]~input_o  = hps_f2h_sdram0_data_writedata[44];

assign \hps_f2h_sdram0_data_writedata[45]~input_o  = hps_f2h_sdram0_data_writedata[45];

assign \hps_f2h_sdram0_data_writedata[46]~input_o  = hps_f2h_sdram0_data_writedata[46];

assign \hps_f2h_sdram0_data_writedata[47]~input_o  = hps_f2h_sdram0_data_writedata[47];

assign \hps_f2h_sdram0_data_writedata[48]~input_o  = hps_f2h_sdram0_data_writedata[48];

assign \hps_f2h_sdram0_data_writedata[49]~input_o  = hps_f2h_sdram0_data_writedata[49];

assign \hps_f2h_sdram0_data_writedata[50]~input_o  = hps_f2h_sdram0_data_writedata[50];

assign \hps_f2h_sdram0_data_writedata[51]~input_o  = hps_f2h_sdram0_data_writedata[51];

assign \hps_f2h_sdram0_data_writedata[52]~input_o  = hps_f2h_sdram0_data_writedata[52];

assign \hps_f2h_sdram0_data_writedata[53]~input_o  = hps_f2h_sdram0_data_writedata[53];

assign \hps_f2h_sdram0_data_writedata[54]~input_o  = hps_f2h_sdram0_data_writedata[54];

assign \hps_f2h_sdram0_data_writedata[55]~input_o  = hps_f2h_sdram0_data_writedata[55];

assign \hps_f2h_sdram0_data_writedata[56]~input_o  = hps_f2h_sdram0_data_writedata[56];

assign \hps_f2h_sdram0_data_writedata[57]~input_o  = hps_f2h_sdram0_data_writedata[57];

assign \hps_f2h_sdram0_data_writedata[58]~input_o  = hps_f2h_sdram0_data_writedata[58];

assign \hps_f2h_sdram0_data_writedata[59]~input_o  = hps_f2h_sdram0_data_writedata[59];

assign \hps_f2h_sdram0_data_writedata[60]~input_o  = hps_f2h_sdram0_data_writedata[60];

assign \hps_f2h_sdram0_data_writedata[61]~input_o  = hps_f2h_sdram0_data_writedata[61];

assign \hps_f2h_sdram0_data_writedata[62]~input_o  = hps_f2h_sdram0_data_writedata[62];

assign \hps_f2h_sdram0_data_writedata[63]~input_o  = hps_f2h_sdram0_data_writedata[63];

assign \hps_f2h_sdram0_data_byteenable[0]~input_o  = hps_f2h_sdram0_data_byteenable[0];

assign \hps_f2h_sdram0_data_byteenable[1]~input_o  = hps_f2h_sdram0_data_byteenable[1];

assign \hps_f2h_sdram0_data_byteenable[2]~input_o  = hps_f2h_sdram0_data_byteenable[2];

assign \hps_f2h_sdram0_data_byteenable[3]~input_o  = hps_f2h_sdram0_data_byteenable[3];

assign \hps_f2h_sdram0_data_byteenable[4]~input_o  = hps_f2h_sdram0_data_byteenable[4];

assign \hps_f2h_sdram0_data_byteenable[5]~input_o  = hps_f2h_sdram0_data_byteenable[5];

assign \hps_f2h_sdram0_data_byteenable[6]~input_o  = hps_f2h_sdram0_data_byteenable[6];

assign \hps_f2h_sdram0_data_byteenable[7]~input_o  = hps_f2h_sdram0_data_byteenable[7];

assign \hps_f2h_sdram0_data_writedata[64]~input_o  = hps_f2h_sdram0_data_writedata[64];

assign \hps_f2h_sdram0_data_writedata[65]~input_o  = hps_f2h_sdram0_data_writedata[65];

assign \hps_f2h_sdram0_data_writedata[66]~input_o  = hps_f2h_sdram0_data_writedata[66];

assign \hps_f2h_sdram0_data_writedata[67]~input_o  = hps_f2h_sdram0_data_writedata[67];

assign \hps_f2h_sdram0_data_writedata[68]~input_o  = hps_f2h_sdram0_data_writedata[68];

assign \hps_f2h_sdram0_data_writedata[69]~input_o  = hps_f2h_sdram0_data_writedata[69];

assign \hps_f2h_sdram0_data_writedata[70]~input_o  = hps_f2h_sdram0_data_writedata[70];

assign \hps_f2h_sdram0_data_writedata[71]~input_o  = hps_f2h_sdram0_data_writedata[71];

assign \hps_f2h_sdram0_data_writedata[72]~input_o  = hps_f2h_sdram0_data_writedata[72];

assign \hps_f2h_sdram0_data_writedata[73]~input_o  = hps_f2h_sdram0_data_writedata[73];

assign \hps_f2h_sdram0_data_writedata[74]~input_o  = hps_f2h_sdram0_data_writedata[74];

assign \hps_f2h_sdram0_data_writedata[75]~input_o  = hps_f2h_sdram0_data_writedata[75];

assign \hps_f2h_sdram0_data_writedata[76]~input_o  = hps_f2h_sdram0_data_writedata[76];

assign \hps_f2h_sdram0_data_writedata[77]~input_o  = hps_f2h_sdram0_data_writedata[77];

assign \hps_f2h_sdram0_data_writedata[78]~input_o  = hps_f2h_sdram0_data_writedata[78];

assign \hps_f2h_sdram0_data_writedata[79]~input_o  = hps_f2h_sdram0_data_writedata[79];

assign \hps_f2h_sdram0_data_writedata[80]~input_o  = hps_f2h_sdram0_data_writedata[80];

assign \hps_f2h_sdram0_data_writedata[81]~input_o  = hps_f2h_sdram0_data_writedata[81];

assign \hps_f2h_sdram0_data_writedata[82]~input_o  = hps_f2h_sdram0_data_writedata[82];

assign \hps_f2h_sdram0_data_writedata[83]~input_o  = hps_f2h_sdram0_data_writedata[83];

assign \hps_f2h_sdram0_data_writedata[84]~input_o  = hps_f2h_sdram0_data_writedata[84];

assign \hps_f2h_sdram0_data_writedata[85]~input_o  = hps_f2h_sdram0_data_writedata[85];

assign \hps_f2h_sdram0_data_writedata[86]~input_o  = hps_f2h_sdram0_data_writedata[86];

assign \hps_f2h_sdram0_data_writedata[87]~input_o  = hps_f2h_sdram0_data_writedata[87];

assign \hps_f2h_sdram0_data_writedata[88]~input_o  = hps_f2h_sdram0_data_writedata[88];

assign \hps_f2h_sdram0_data_writedata[89]~input_o  = hps_f2h_sdram0_data_writedata[89];

assign \hps_f2h_sdram0_data_writedata[90]~input_o  = hps_f2h_sdram0_data_writedata[90];

assign \hps_f2h_sdram0_data_writedata[91]~input_o  = hps_f2h_sdram0_data_writedata[91];

assign \hps_f2h_sdram0_data_writedata[92]~input_o  = hps_f2h_sdram0_data_writedata[92];

assign \hps_f2h_sdram0_data_writedata[93]~input_o  = hps_f2h_sdram0_data_writedata[93];

assign \hps_f2h_sdram0_data_writedata[94]~input_o  = hps_f2h_sdram0_data_writedata[94];

assign \hps_f2h_sdram0_data_writedata[95]~input_o  = hps_f2h_sdram0_data_writedata[95];

assign \hps_f2h_sdram0_data_writedata[96]~input_o  = hps_f2h_sdram0_data_writedata[96];

assign \hps_f2h_sdram0_data_writedata[97]~input_o  = hps_f2h_sdram0_data_writedata[97];

assign \hps_f2h_sdram0_data_writedata[98]~input_o  = hps_f2h_sdram0_data_writedata[98];

assign \hps_f2h_sdram0_data_writedata[99]~input_o  = hps_f2h_sdram0_data_writedata[99];

assign \hps_f2h_sdram0_data_writedata[100]~input_o  = hps_f2h_sdram0_data_writedata[100];

assign \hps_f2h_sdram0_data_writedata[101]~input_o  = hps_f2h_sdram0_data_writedata[101];

assign \hps_f2h_sdram0_data_writedata[102]~input_o  = hps_f2h_sdram0_data_writedata[102];

assign \hps_f2h_sdram0_data_writedata[103]~input_o  = hps_f2h_sdram0_data_writedata[103];

assign \hps_f2h_sdram0_data_writedata[104]~input_o  = hps_f2h_sdram0_data_writedata[104];

assign \hps_f2h_sdram0_data_writedata[105]~input_o  = hps_f2h_sdram0_data_writedata[105];

assign \hps_f2h_sdram0_data_writedata[106]~input_o  = hps_f2h_sdram0_data_writedata[106];

assign \hps_f2h_sdram0_data_writedata[107]~input_o  = hps_f2h_sdram0_data_writedata[107];

assign \hps_f2h_sdram0_data_writedata[108]~input_o  = hps_f2h_sdram0_data_writedata[108];

assign \hps_f2h_sdram0_data_writedata[109]~input_o  = hps_f2h_sdram0_data_writedata[109];

assign \hps_f2h_sdram0_data_writedata[110]~input_o  = hps_f2h_sdram0_data_writedata[110];

assign \hps_f2h_sdram0_data_writedata[111]~input_o  = hps_f2h_sdram0_data_writedata[111];

assign \hps_f2h_sdram0_data_writedata[112]~input_o  = hps_f2h_sdram0_data_writedata[112];

assign \hps_f2h_sdram0_data_writedata[113]~input_o  = hps_f2h_sdram0_data_writedata[113];

assign \hps_f2h_sdram0_data_writedata[114]~input_o  = hps_f2h_sdram0_data_writedata[114];

assign \hps_f2h_sdram0_data_writedata[115]~input_o  = hps_f2h_sdram0_data_writedata[115];

assign \hps_f2h_sdram0_data_writedata[116]~input_o  = hps_f2h_sdram0_data_writedata[116];

assign \hps_f2h_sdram0_data_writedata[117]~input_o  = hps_f2h_sdram0_data_writedata[117];

assign \hps_f2h_sdram0_data_writedata[118]~input_o  = hps_f2h_sdram0_data_writedata[118];

assign \hps_f2h_sdram0_data_writedata[119]~input_o  = hps_f2h_sdram0_data_writedata[119];

assign \hps_f2h_sdram0_data_writedata[120]~input_o  = hps_f2h_sdram0_data_writedata[120];

assign \hps_f2h_sdram0_data_writedata[121]~input_o  = hps_f2h_sdram0_data_writedata[121];

assign \hps_f2h_sdram0_data_writedata[122]~input_o  = hps_f2h_sdram0_data_writedata[122];

assign \hps_f2h_sdram0_data_writedata[123]~input_o  = hps_f2h_sdram0_data_writedata[123];

assign \hps_f2h_sdram0_data_writedata[124]~input_o  = hps_f2h_sdram0_data_writedata[124];

assign \hps_f2h_sdram0_data_writedata[125]~input_o  = hps_f2h_sdram0_data_writedata[125];

assign \hps_f2h_sdram0_data_writedata[126]~input_o  = hps_f2h_sdram0_data_writedata[126];

assign \hps_f2h_sdram0_data_writedata[127]~input_o  = hps_f2h_sdram0_data_writedata[127];

assign \hps_f2h_sdram0_data_byteenable[8]~input_o  = hps_f2h_sdram0_data_byteenable[8];

assign \hps_f2h_sdram0_data_byteenable[9]~input_o  = hps_f2h_sdram0_data_byteenable[9];

assign \hps_f2h_sdram0_data_byteenable[10]~input_o  = hps_f2h_sdram0_data_byteenable[10];

assign \hps_f2h_sdram0_data_byteenable[11]~input_o  = hps_f2h_sdram0_data_byteenable[11];

assign \hps_f2h_sdram0_data_byteenable[12]~input_o  = hps_f2h_sdram0_data_byteenable[12];

assign \hps_f2h_sdram0_data_byteenable[13]~input_o  = hps_f2h_sdram0_data_byteenable[13];

assign \hps_f2h_sdram0_data_byteenable[14]~input_o  = hps_f2h_sdram0_data_byteenable[14];

assign \hps_f2h_sdram0_data_byteenable[15]~input_o  = hps_f2h_sdram0_data_byteenable[15];

assign \hps_f2h_sdram0_data_writedata[128]~input_o  = hps_f2h_sdram0_data_writedata[128];

assign \hps_f2h_sdram0_data_writedata[129]~input_o  = hps_f2h_sdram0_data_writedata[129];

assign \hps_f2h_sdram0_data_writedata[130]~input_o  = hps_f2h_sdram0_data_writedata[130];

assign \hps_f2h_sdram0_data_writedata[131]~input_o  = hps_f2h_sdram0_data_writedata[131];

assign \hps_f2h_sdram0_data_writedata[132]~input_o  = hps_f2h_sdram0_data_writedata[132];

assign \hps_f2h_sdram0_data_writedata[133]~input_o  = hps_f2h_sdram0_data_writedata[133];

assign \hps_f2h_sdram0_data_writedata[134]~input_o  = hps_f2h_sdram0_data_writedata[134];

assign \hps_f2h_sdram0_data_writedata[135]~input_o  = hps_f2h_sdram0_data_writedata[135];

assign \hps_f2h_sdram0_data_writedata[136]~input_o  = hps_f2h_sdram0_data_writedata[136];

assign \hps_f2h_sdram0_data_writedata[137]~input_o  = hps_f2h_sdram0_data_writedata[137];

assign \hps_f2h_sdram0_data_writedata[138]~input_o  = hps_f2h_sdram0_data_writedata[138];

assign \hps_f2h_sdram0_data_writedata[139]~input_o  = hps_f2h_sdram0_data_writedata[139];

assign \hps_f2h_sdram0_data_writedata[140]~input_o  = hps_f2h_sdram0_data_writedata[140];

assign \hps_f2h_sdram0_data_writedata[141]~input_o  = hps_f2h_sdram0_data_writedata[141];

assign \hps_f2h_sdram0_data_writedata[142]~input_o  = hps_f2h_sdram0_data_writedata[142];

assign \hps_f2h_sdram0_data_writedata[143]~input_o  = hps_f2h_sdram0_data_writedata[143];

assign \hps_f2h_sdram0_data_writedata[144]~input_o  = hps_f2h_sdram0_data_writedata[144];

assign \hps_f2h_sdram0_data_writedata[145]~input_o  = hps_f2h_sdram0_data_writedata[145];

assign \hps_f2h_sdram0_data_writedata[146]~input_o  = hps_f2h_sdram0_data_writedata[146];

assign \hps_f2h_sdram0_data_writedata[147]~input_o  = hps_f2h_sdram0_data_writedata[147];

assign \hps_f2h_sdram0_data_writedata[148]~input_o  = hps_f2h_sdram0_data_writedata[148];

assign \hps_f2h_sdram0_data_writedata[149]~input_o  = hps_f2h_sdram0_data_writedata[149];

assign \hps_f2h_sdram0_data_writedata[150]~input_o  = hps_f2h_sdram0_data_writedata[150];

assign \hps_f2h_sdram0_data_writedata[151]~input_o  = hps_f2h_sdram0_data_writedata[151];

assign \hps_f2h_sdram0_data_writedata[152]~input_o  = hps_f2h_sdram0_data_writedata[152];

assign \hps_f2h_sdram0_data_writedata[153]~input_o  = hps_f2h_sdram0_data_writedata[153];

assign \hps_f2h_sdram0_data_writedata[154]~input_o  = hps_f2h_sdram0_data_writedata[154];

assign \hps_f2h_sdram0_data_writedata[155]~input_o  = hps_f2h_sdram0_data_writedata[155];

assign \hps_f2h_sdram0_data_writedata[156]~input_o  = hps_f2h_sdram0_data_writedata[156];

assign \hps_f2h_sdram0_data_writedata[157]~input_o  = hps_f2h_sdram0_data_writedata[157];

assign \hps_f2h_sdram0_data_writedata[158]~input_o  = hps_f2h_sdram0_data_writedata[158];

assign \hps_f2h_sdram0_data_writedata[159]~input_o  = hps_f2h_sdram0_data_writedata[159];

assign \hps_f2h_sdram0_data_writedata[160]~input_o  = hps_f2h_sdram0_data_writedata[160];

assign \hps_f2h_sdram0_data_writedata[161]~input_o  = hps_f2h_sdram0_data_writedata[161];

assign \hps_f2h_sdram0_data_writedata[162]~input_o  = hps_f2h_sdram0_data_writedata[162];

assign \hps_f2h_sdram0_data_writedata[163]~input_o  = hps_f2h_sdram0_data_writedata[163];

assign \hps_f2h_sdram0_data_writedata[164]~input_o  = hps_f2h_sdram0_data_writedata[164];

assign \hps_f2h_sdram0_data_writedata[165]~input_o  = hps_f2h_sdram0_data_writedata[165];

assign \hps_f2h_sdram0_data_writedata[166]~input_o  = hps_f2h_sdram0_data_writedata[166];

assign \hps_f2h_sdram0_data_writedata[167]~input_o  = hps_f2h_sdram0_data_writedata[167];

assign \hps_f2h_sdram0_data_writedata[168]~input_o  = hps_f2h_sdram0_data_writedata[168];

assign \hps_f2h_sdram0_data_writedata[169]~input_o  = hps_f2h_sdram0_data_writedata[169];

assign \hps_f2h_sdram0_data_writedata[170]~input_o  = hps_f2h_sdram0_data_writedata[170];

assign \hps_f2h_sdram0_data_writedata[171]~input_o  = hps_f2h_sdram0_data_writedata[171];

assign \hps_f2h_sdram0_data_writedata[172]~input_o  = hps_f2h_sdram0_data_writedata[172];

assign \hps_f2h_sdram0_data_writedata[173]~input_o  = hps_f2h_sdram0_data_writedata[173];

assign \hps_f2h_sdram0_data_writedata[174]~input_o  = hps_f2h_sdram0_data_writedata[174];

assign \hps_f2h_sdram0_data_writedata[175]~input_o  = hps_f2h_sdram0_data_writedata[175];

assign \hps_f2h_sdram0_data_writedata[176]~input_o  = hps_f2h_sdram0_data_writedata[176];

assign \hps_f2h_sdram0_data_writedata[177]~input_o  = hps_f2h_sdram0_data_writedata[177];

assign \hps_f2h_sdram0_data_writedata[178]~input_o  = hps_f2h_sdram0_data_writedata[178];

assign \hps_f2h_sdram0_data_writedata[179]~input_o  = hps_f2h_sdram0_data_writedata[179];

assign \hps_f2h_sdram0_data_writedata[180]~input_o  = hps_f2h_sdram0_data_writedata[180];

assign \hps_f2h_sdram0_data_writedata[181]~input_o  = hps_f2h_sdram0_data_writedata[181];

assign \hps_f2h_sdram0_data_writedata[182]~input_o  = hps_f2h_sdram0_data_writedata[182];

assign \hps_f2h_sdram0_data_writedata[183]~input_o  = hps_f2h_sdram0_data_writedata[183];

assign \hps_f2h_sdram0_data_writedata[184]~input_o  = hps_f2h_sdram0_data_writedata[184];

assign \hps_f2h_sdram0_data_writedata[185]~input_o  = hps_f2h_sdram0_data_writedata[185];

assign \hps_f2h_sdram0_data_writedata[186]~input_o  = hps_f2h_sdram0_data_writedata[186];

assign \hps_f2h_sdram0_data_writedata[187]~input_o  = hps_f2h_sdram0_data_writedata[187];

assign \hps_f2h_sdram0_data_writedata[188]~input_o  = hps_f2h_sdram0_data_writedata[188];

assign \hps_f2h_sdram0_data_writedata[189]~input_o  = hps_f2h_sdram0_data_writedata[189];

assign \hps_f2h_sdram0_data_writedata[190]~input_o  = hps_f2h_sdram0_data_writedata[190];

assign \hps_f2h_sdram0_data_writedata[191]~input_o  = hps_f2h_sdram0_data_writedata[191];

assign \hps_f2h_sdram0_data_byteenable[16]~input_o  = hps_f2h_sdram0_data_byteenable[16];

assign \hps_f2h_sdram0_data_byteenable[17]~input_o  = hps_f2h_sdram0_data_byteenable[17];

assign \hps_f2h_sdram0_data_byteenable[18]~input_o  = hps_f2h_sdram0_data_byteenable[18];

assign \hps_f2h_sdram0_data_byteenable[19]~input_o  = hps_f2h_sdram0_data_byteenable[19];

assign \hps_f2h_sdram0_data_byteenable[20]~input_o  = hps_f2h_sdram0_data_byteenable[20];

assign \hps_f2h_sdram0_data_byteenable[21]~input_o  = hps_f2h_sdram0_data_byteenable[21];

assign \hps_f2h_sdram0_data_byteenable[22]~input_o  = hps_f2h_sdram0_data_byteenable[22];

assign \hps_f2h_sdram0_data_byteenable[23]~input_o  = hps_f2h_sdram0_data_byteenable[23];

assign \hps_f2h_sdram0_data_writedata[192]~input_o  = hps_f2h_sdram0_data_writedata[192];

assign \hps_f2h_sdram0_data_writedata[193]~input_o  = hps_f2h_sdram0_data_writedata[193];

assign \hps_f2h_sdram0_data_writedata[194]~input_o  = hps_f2h_sdram0_data_writedata[194];

assign \hps_f2h_sdram0_data_writedata[195]~input_o  = hps_f2h_sdram0_data_writedata[195];

assign \hps_f2h_sdram0_data_writedata[196]~input_o  = hps_f2h_sdram0_data_writedata[196];

assign \hps_f2h_sdram0_data_writedata[197]~input_o  = hps_f2h_sdram0_data_writedata[197];

assign \hps_f2h_sdram0_data_writedata[198]~input_o  = hps_f2h_sdram0_data_writedata[198];

assign \hps_f2h_sdram0_data_writedata[199]~input_o  = hps_f2h_sdram0_data_writedata[199];

assign \hps_f2h_sdram0_data_writedata[200]~input_o  = hps_f2h_sdram0_data_writedata[200];

assign \hps_f2h_sdram0_data_writedata[201]~input_o  = hps_f2h_sdram0_data_writedata[201];

assign \hps_f2h_sdram0_data_writedata[202]~input_o  = hps_f2h_sdram0_data_writedata[202];

assign \hps_f2h_sdram0_data_writedata[203]~input_o  = hps_f2h_sdram0_data_writedata[203];

assign \hps_f2h_sdram0_data_writedata[204]~input_o  = hps_f2h_sdram0_data_writedata[204];

assign \hps_f2h_sdram0_data_writedata[205]~input_o  = hps_f2h_sdram0_data_writedata[205];

assign \hps_f2h_sdram0_data_writedata[206]~input_o  = hps_f2h_sdram0_data_writedata[206];

assign \hps_f2h_sdram0_data_writedata[207]~input_o  = hps_f2h_sdram0_data_writedata[207];

assign \hps_f2h_sdram0_data_writedata[208]~input_o  = hps_f2h_sdram0_data_writedata[208];

assign \hps_f2h_sdram0_data_writedata[209]~input_o  = hps_f2h_sdram0_data_writedata[209];

assign \hps_f2h_sdram0_data_writedata[210]~input_o  = hps_f2h_sdram0_data_writedata[210];

assign \hps_f2h_sdram0_data_writedata[211]~input_o  = hps_f2h_sdram0_data_writedata[211];

assign \hps_f2h_sdram0_data_writedata[212]~input_o  = hps_f2h_sdram0_data_writedata[212];

assign \hps_f2h_sdram0_data_writedata[213]~input_o  = hps_f2h_sdram0_data_writedata[213];

assign \hps_f2h_sdram0_data_writedata[214]~input_o  = hps_f2h_sdram0_data_writedata[214];

assign \hps_f2h_sdram0_data_writedata[215]~input_o  = hps_f2h_sdram0_data_writedata[215];

assign \hps_f2h_sdram0_data_writedata[216]~input_o  = hps_f2h_sdram0_data_writedata[216];

assign \hps_f2h_sdram0_data_writedata[217]~input_o  = hps_f2h_sdram0_data_writedata[217];

assign \hps_f2h_sdram0_data_writedata[218]~input_o  = hps_f2h_sdram0_data_writedata[218];

assign \hps_f2h_sdram0_data_writedata[219]~input_o  = hps_f2h_sdram0_data_writedata[219];

assign \hps_f2h_sdram0_data_writedata[220]~input_o  = hps_f2h_sdram0_data_writedata[220];

assign \hps_f2h_sdram0_data_writedata[221]~input_o  = hps_f2h_sdram0_data_writedata[221];

assign \hps_f2h_sdram0_data_writedata[222]~input_o  = hps_f2h_sdram0_data_writedata[222];

assign \hps_f2h_sdram0_data_writedata[223]~input_o  = hps_f2h_sdram0_data_writedata[223];

assign \hps_f2h_sdram0_data_writedata[224]~input_o  = hps_f2h_sdram0_data_writedata[224];

assign \hps_f2h_sdram0_data_writedata[225]~input_o  = hps_f2h_sdram0_data_writedata[225];

assign \hps_f2h_sdram0_data_writedata[226]~input_o  = hps_f2h_sdram0_data_writedata[226];

assign \hps_f2h_sdram0_data_writedata[227]~input_o  = hps_f2h_sdram0_data_writedata[227];

assign \hps_f2h_sdram0_data_writedata[228]~input_o  = hps_f2h_sdram0_data_writedata[228];

assign \hps_f2h_sdram0_data_writedata[229]~input_o  = hps_f2h_sdram0_data_writedata[229];

assign \hps_f2h_sdram0_data_writedata[230]~input_o  = hps_f2h_sdram0_data_writedata[230];

assign \hps_f2h_sdram0_data_writedata[231]~input_o  = hps_f2h_sdram0_data_writedata[231];

assign \hps_f2h_sdram0_data_writedata[232]~input_o  = hps_f2h_sdram0_data_writedata[232];

assign \hps_f2h_sdram0_data_writedata[233]~input_o  = hps_f2h_sdram0_data_writedata[233];

assign \hps_f2h_sdram0_data_writedata[234]~input_o  = hps_f2h_sdram0_data_writedata[234];

assign \hps_f2h_sdram0_data_writedata[235]~input_o  = hps_f2h_sdram0_data_writedata[235];

assign \hps_f2h_sdram0_data_writedata[236]~input_o  = hps_f2h_sdram0_data_writedata[236];

assign \hps_f2h_sdram0_data_writedata[237]~input_o  = hps_f2h_sdram0_data_writedata[237];

assign \hps_f2h_sdram0_data_writedata[238]~input_o  = hps_f2h_sdram0_data_writedata[238];

assign \hps_f2h_sdram0_data_writedata[239]~input_o  = hps_f2h_sdram0_data_writedata[239];

assign \hps_f2h_sdram0_data_writedata[240]~input_o  = hps_f2h_sdram0_data_writedata[240];

assign \hps_f2h_sdram0_data_writedata[241]~input_o  = hps_f2h_sdram0_data_writedata[241];

assign \hps_f2h_sdram0_data_writedata[242]~input_o  = hps_f2h_sdram0_data_writedata[242];

assign \hps_f2h_sdram0_data_writedata[243]~input_o  = hps_f2h_sdram0_data_writedata[243];

assign \hps_f2h_sdram0_data_writedata[244]~input_o  = hps_f2h_sdram0_data_writedata[244];

assign \hps_f2h_sdram0_data_writedata[245]~input_o  = hps_f2h_sdram0_data_writedata[245];

assign \hps_f2h_sdram0_data_writedata[246]~input_o  = hps_f2h_sdram0_data_writedata[246];

assign \hps_f2h_sdram0_data_writedata[247]~input_o  = hps_f2h_sdram0_data_writedata[247];

assign \hps_f2h_sdram0_data_writedata[248]~input_o  = hps_f2h_sdram0_data_writedata[248];

assign \hps_f2h_sdram0_data_writedata[249]~input_o  = hps_f2h_sdram0_data_writedata[249];

assign \hps_f2h_sdram0_data_writedata[250]~input_o  = hps_f2h_sdram0_data_writedata[250];

assign \hps_f2h_sdram0_data_writedata[251]~input_o  = hps_f2h_sdram0_data_writedata[251];

assign \hps_f2h_sdram0_data_writedata[252]~input_o  = hps_f2h_sdram0_data_writedata[252];

assign \hps_f2h_sdram0_data_writedata[253]~input_o  = hps_f2h_sdram0_data_writedata[253];

assign \hps_f2h_sdram0_data_writedata[254]~input_o  = hps_f2h_sdram0_data_writedata[254];

assign \hps_f2h_sdram0_data_writedata[255]~input_o  = hps_f2h_sdram0_data_writedata[255];

assign \hps_f2h_sdram0_data_byteenable[24]~input_o  = hps_f2h_sdram0_data_byteenable[24];

assign \hps_f2h_sdram0_data_byteenable[25]~input_o  = hps_f2h_sdram0_data_byteenable[25];

assign \hps_f2h_sdram0_data_byteenable[26]~input_o  = hps_f2h_sdram0_data_byteenable[26];

assign \hps_f2h_sdram0_data_byteenable[27]~input_o  = hps_f2h_sdram0_data_byteenable[27];

assign \hps_f2h_sdram0_data_byteenable[28]~input_o  = hps_f2h_sdram0_data_byteenable[28];

assign \hps_f2h_sdram0_data_byteenable[29]~input_o  = hps_f2h_sdram0_data_byteenable[29];

assign \hps_f2h_sdram0_data_byteenable[30]~input_o  = hps_f2h_sdram0_data_byteenable[30];

assign \hps_f2h_sdram0_data_byteenable[31]~input_o  = hps_f2h_sdram0_data_byteenable[31];

assign \reset_reset_n~input_o  = reset_reset_n;

assign \state_in_export[0]~input_o  = state_in_export[0];

assign \switches_in_export[0]~input_o  = switches_in_export[0];

assign \state_in_export[1]~input_o  = state_in_export[1];

assign \switches_in_export[1]~input_o  = switches_in_export[1];

assign \state_in_export[2]~input_o  = state_in_export[2];

assign \switches_in_export[2]~input_o  = switches_in_export[2];

assign \state_in_export[3]~input_o  = state_in_export[3];

assign \switches_in_export[3]~input_o  = switches_in_export[3];

assign \state_in_export[4]~input_o  = state_in_export[4];

assign \switches_in_export[4]~input_o  = switches_in_export[4];

assign \state_in_export[5]~input_o  = state_in_export[5];

assign \switches_in_export[5]~input_o  = switches_in_export[5];

assign \state_in_export[6]~input_o  = state_in_export[6];

assign \switches_in_export[6]~input_o  = switches_in_export[6];

assign \state_in_export[7]~input_o  = state_in_export[7];

assign \switches_in_export[7]~input_o  = switches_in_export[7];

assign \state_in_export[8]~input_o  = state_in_export[8];

assign \switches_in_export[8]~input_o  = switches_in_export[8];

assign \state_in_export[9]~input_o  = state_in_export[9];

assign \switches_in_export[9]~input_o  = switches_in_export[9];

assign \state_in_export[10]~input_o  = state_in_export[10];

assign \state_in_export[11]~input_o  = state_in_export[11];

assign \state_in_export[12]~input_o  = state_in_export[12];

assign \state_in_export[13]~input_o  = state_in_export[13];

assign \state_in_export[14]~input_o  = state_in_export[14];

assign \state_in_export[15]~input_o  = state_in_export[15];

assign \state_in_export[16]~input_o  = state_in_export[16];

assign \state_in_export[17]~input_o  = state_in_export[17];

assign \state_in_export[18]~input_o  = state_in_export[18];

assign \state_in_export[19]~input_o  = state_in_export[19];

assign \state_in_export[20]~input_o  = state_in_export[20];

assign \state_in_export[21]~input_o  = state_in_export[21];

assign \state_in_export[22]~input_o  = state_in_export[22];

assign \state_in_export[23]~input_o  = state_in_export[23];

assign \state_in_export[24]~input_o  = state_in_export[24];

assign \state_in_export[25]~input_o  = state_in_export[25];

assign \state_in_export[26]~input_o  = state_in_export[26];

assign \state_in_export[27]~input_o  = state_in_export[27];

assign \state_in_export[28]~input_o  = state_in_export[28];

assign \state_in_export[29]~input_o  = state_in_export[29];

assign \state_in_export[30]~input_o  = state_in_export[30];

assign \state_in_export[31]~input_o  = state_in_export[31];

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[3]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[2]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[1]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].delayed_data_out ),
	.oe(vcc),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dm[0]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|extra_output_pad_gen[0].obuf_1 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_obar[0] ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oebout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck_n),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obuf_ba_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_o[0] ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|wire_pseudo_diffa_oeout[0] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(memory_mem_ck),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|clock_gen[0].uclk_generator|obufa_0 .shift_series_termination_control = "false";

assign base_addr_ddr_out_export[0] = \base_address_ddr|data_out[0]~q ;

assign base_addr_ddr_out_export[1] = \base_address_ddr|data_out[1]~q ;

assign base_addr_ddr_out_export[2] = \base_address_ddr|data_out[2]~q ;

assign base_addr_ddr_out_export[3] = \base_address_ddr|data_out[3]~q ;

assign base_addr_ddr_out_export[4] = \base_address_ddr|data_out[4]~q ;

assign base_addr_ddr_out_export[5] = \base_address_ddr|data_out[5]~q ;

assign base_addr_ddr_out_export[6] = \base_address_ddr|data_out[6]~q ;

assign base_addr_ddr_out_export[7] = \base_address_ddr|data_out[7]~q ;

assign base_addr_ddr_out_export[8] = \base_address_ddr|data_out[8]~q ;

assign base_addr_ddr_out_export[9] = \base_address_ddr|data_out[9]~q ;

assign base_addr_ddr_out_export[10] = \base_address_ddr|data_out[10]~q ;

assign base_addr_ddr_out_export[11] = \base_address_ddr|data_out[11]~q ;

assign base_addr_ddr_out_export[12] = \base_address_ddr|data_out[12]~q ;

assign base_addr_ddr_out_export[13] = \base_address_ddr|data_out[13]~q ;

assign base_addr_ddr_out_export[14] = \base_address_ddr|data_out[14]~q ;

assign base_addr_ddr_out_export[15] = \base_address_ddr|data_out[15]~q ;

assign base_addr_ddr_out_export[16] = \base_address_ddr|data_out[16]~q ;

assign base_addr_ddr_out_export[17] = \base_address_ddr|data_out[17]~q ;

assign base_addr_ddr_out_export[18] = \base_address_ddr|data_out[18]~q ;

assign base_addr_ddr_out_export[19] = \base_address_ddr|data_out[19]~q ;

assign base_addr_ddr_out_export[20] = \base_address_ddr|data_out[20]~q ;

assign base_addr_ddr_out_export[21] = \base_address_ddr|data_out[21]~q ;

assign base_addr_ddr_out_export[22] = \base_address_ddr|data_out[22]~q ;

assign base_addr_ddr_out_export[23] = \base_address_ddr|data_out[23]~q ;

assign base_addr_ddr_out_export[24] = \base_address_ddr|data_out[24]~q ;

assign base_addr_ddr_out_export[25] = \base_address_ddr|data_out[25]~q ;

assign base_addr_ddr_out_export[26] = \base_address_ddr|data_out[26]~q ;

assign base_addr_ddr_out_export[27] = \base_address_ddr|data_out[27]~q ;

assign base_addr_ddr_out_export[28] = \base_address_ddr|data_out[28]~q ;

assign base_addr_ddr_out_export[29] = \base_address_ddr|data_out[29]~q ;

assign base_addr_ddr_out_export[30] = \base_address_ddr|data_out[30]~q ;

assign base_addr_ddr_out_export[31] = \base_address_ddr|data_out[31]~q ;

assign control_out_export[0] = \control|data_out[0]~q ;

assign control_out_export[1] = \control|data_out[1]~q ;

assign control_out_export[2] = \control|data_out[2]~q ;

assign control_out_export[3] = \control|data_out[3]~q ;

assign control_out_export[4] = \control|data_out[4]~q ;

assign control_out_export[5] = \control|data_out[5]~q ;

assign control_out_export[6] = \control|data_out[6]~q ;

assign control_out_export[7] = \control|data_out[7]~q ;

assign control_out_export[8] = \control|data_out[8]~q ;

assign control_out_export[9] = \control|data_out[9]~q ;

assign control_out_export[10] = \control|data_out[10]~q ;

assign control_out_export[11] = \control|data_out[11]~q ;

assign control_out_export[12] = \control|data_out[12]~q ;

assign control_out_export[13] = \control|data_out[13]~q ;

assign control_out_export[14] = \control|data_out[14]~q ;

assign control_out_export[15] = \control|data_out[15]~q ;

assign control_out_export[16] = \control|data_out[16]~q ;

assign control_out_export[17] = \control|data_out[17]~q ;

assign control_out_export[18] = \control|data_out[18]~q ;

assign control_out_export[19] = \control|data_out[19]~q ;

assign control_out_export[20] = \control|data_out[20]~q ;

assign control_out_export[21] = \control|data_out[21]~q ;

assign control_out_export[22] = \control|data_out[22]~q ;

assign control_out_export[23] = \control|data_out[23]~q ;

assign control_out_export[24] = \control|data_out[24]~q ;

assign control_out_export[25] = \control|data_out[25]~q ;

assign control_out_export[26] = \control|data_out[26]~q ;

assign control_out_export[27] = \control|data_out[27]~q ;

assign control_out_export[28] = \control|data_out[28]~q ;

assign control_out_export[29] = \control|data_out[29]~q ;

assign control_out_export[30] = \control|data_out[30]~q ;

assign control_out_export[31] = \control|data_out[31]~q ;

assign hps_f2h_sdram0_data_waitrequest = ~ \hps|fpga_interfaces|intermediate[1] ;

assign hps_f2h_sdram0_data_readdata[0] = \hps|fpga_interfaces|f2h_sdram0_READDATA[0] ;

assign hps_f2h_sdram0_data_readdata[1] = \hps|fpga_interfaces|f2h_sdram0_READDATA[1] ;

assign hps_f2h_sdram0_data_readdata[2] = \hps|fpga_interfaces|f2h_sdram0_READDATA[2] ;

assign hps_f2h_sdram0_data_readdata[3] = \hps|fpga_interfaces|f2h_sdram0_READDATA[3] ;

assign hps_f2h_sdram0_data_readdata[4] = \hps|fpga_interfaces|f2h_sdram0_READDATA[4] ;

assign hps_f2h_sdram0_data_readdata[5] = \hps|fpga_interfaces|f2h_sdram0_READDATA[5] ;

assign hps_f2h_sdram0_data_readdata[6] = \hps|fpga_interfaces|f2h_sdram0_READDATA[6] ;

assign hps_f2h_sdram0_data_readdata[7] = \hps|fpga_interfaces|f2h_sdram0_READDATA[7] ;

assign hps_f2h_sdram0_data_readdata[8] = \hps|fpga_interfaces|f2h_sdram0_READDATA[8] ;

assign hps_f2h_sdram0_data_readdata[9] = \hps|fpga_interfaces|f2h_sdram0_READDATA[9] ;

assign hps_f2h_sdram0_data_readdata[10] = \hps|fpga_interfaces|f2h_sdram0_READDATA[10] ;

assign hps_f2h_sdram0_data_readdata[11] = \hps|fpga_interfaces|f2h_sdram0_READDATA[11] ;

assign hps_f2h_sdram0_data_readdata[12] = \hps|fpga_interfaces|f2h_sdram0_READDATA[12] ;

assign hps_f2h_sdram0_data_readdata[13] = \hps|fpga_interfaces|f2h_sdram0_READDATA[13] ;

assign hps_f2h_sdram0_data_readdata[14] = \hps|fpga_interfaces|f2h_sdram0_READDATA[14] ;

assign hps_f2h_sdram0_data_readdata[15] = \hps|fpga_interfaces|f2h_sdram0_READDATA[15] ;

assign hps_f2h_sdram0_data_readdata[16] = \hps|fpga_interfaces|f2h_sdram0_READDATA[16] ;

assign hps_f2h_sdram0_data_readdata[17] = \hps|fpga_interfaces|f2h_sdram0_READDATA[17] ;

assign hps_f2h_sdram0_data_readdata[18] = \hps|fpga_interfaces|f2h_sdram0_READDATA[18] ;

assign hps_f2h_sdram0_data_readdata[19] = \hps|fpga_interfaces|f2h_sdram0_READDATA[19] ;

assign hps_f2h_sdram0_data_readdata[20] = \hps|fpga_interfaces|f2h_sdram0_READDATA[20] ;

assign hps_f2h_sdram0_data_readdata[21] = \hps|fpga_interfaces|f2h_sdram0_READDATA[21] ;

assign hps_f2h_sdram0_data_readdata[22] = \hps|fpga_interfaces|f2h_sdram0_READDATA[22] ;

assign hps_f2h_sdram0_data_readdata[23] = \hps|fpga_interfaces|f2h_sdram0_READDATA[23] ;

assign hps_f2h_sdram0_data_readdata[24] = \hps|fpga_interfaces|f2h_sdram0_READDATA[24] ;

assign hps_f2h_sdram0_data_readdata[25] = \hps|fpga_interfaces|f2h_sdram0_READDATA[25] ;

assign hps_f2h_sdram0_data_readdata[26] = \hps|fpga_interfaces|f2h_sdram0_READDATA[26] ;

assign hps_f2h_sdram0_data_readdata[27] = \hps|fpga_interfaces|f2h_sdram0_READDATA[27] ;

assign hps_f2h_sdram0_data_readdata[28] = \hps|fpga_interfaces|f2h_sdram0_READDATA[28] ;

assign hps_f2h_sdram0_data_readdata[29] = \hps|fpga_interfaces|f2h_sdram0_READDATA[29] ;

assign hps_f2h_sdram0_data_readdata[30] = \hps|fpga_interfaces|f2h_sdram0_READDATA[30] ;

assign hps_f2h_sdram0_data_readdata[31] = \hps|fpga_interfaces|f2h_sdram0_READDATA[31] ;

assign hps_f2h_sdram0_data_readdata[32] = \hps|fpga_interfaces|f2h_sdram0_READDATA[32] ;

assign hps_f2h_sdram0_data_readdata[33] = \hps|fpga_interfaces|f2h_sdram0_READDATA[33] ;

assign hps_f2h_sdram0_data_readdata[34] = \hps|fpga_interfaces|f2h_sdram0_READDATA[34] ;

assign hps_f2h_sdram0_data_readdata[35] = \hps|fpga_interfaces|f2h_sdram0_READDATA[35] ;

assign hps_f2h_sdram0_data_readdata[36] = \hps|fpga_interfaces|f2h_sdram0_READDATA[36] ;

assign hps_f2h_sdram0_data_readdata[37] = \hps|fpga_interfaces|f2h_sdram0_READDATA[37] ;

assign hps_f2h_sdram0_data_readdata[38] = \hps|fpga_interfaces|f2h_sdram0_READDATA[38] ;

assign hps_f2h_sdram0_data_readdata[39] = \hps|fpga_interfaces|f2h_sdram0_READDATA[39] ;

assign hps_f2h_sdram0_data_readdata[40] = \hps|fpga_interfaces|f2h_sdram0_READDATA[40] ;

assign hps_f2h_sdram0_data_readdata[41] = \hps|fpga_interfaces|f2h_sdram0_READDATA[41] ;

assign hps_f2h_sdram0_data_readdata[42] = \hps|fpga_interfaces|f2h_sdram0_READDATA[42] ;

assign hps_f2h_sdram0_data_readdata[43] = \hps|fpga_interfaces|f2h_sdram0_READDATA[43] ;

assign hps_f2h_sdram0_data_readdata[44] = \hps|fpga_interfaces|f2h_sdram0_READDATA[44] ;

assign hps_f2h_sdram0_data_readdata[45] = \hps|fpga_interfaces|f2h_sdram0_READDATA[45] ;

assign hps_f2h_sdram0_data_readdata[46] = \hps|fpga_interfaces|f2h_sdram0_READDATA[46] ;

assign hps_f2h_sdram0_data_readdata[47] = \hps|fpga_interfaces|f2h_sdram0_READDATA[47] ;

assign hps_f2h_sdram0_data_readdata[48] = \hps|fpga_interfaces|f2h_sdram0_READDATA[48] ;

assign hps_f2h_sdram0_data_readdata[49] = \hps|fpga_interfaces|f2h_sdram0_READDATA[49] ;

assign hps_f2h_sdram0_data_readdata[50] = \hps|fpga_interfaces|f2h_sdram0_READDATA[50] ;

assign hps_f2h_sdram0_data_readdata[51] = \hps|fpga_interfaces|f2h_sdram0_READDATA[51] ;

assign hps_f2h_sdram0_data_readdata[52] = \hps|fpga_interfaces|f2h_sdram0_READDATA[52] ;

assign hps_f2h_sdram0_data_readdata[53] = \hps|fpga_interfaces|f2h_sdram0_READDATA[53] ;

assign hps_f2h_sdram0_data_readdata[54] = \hps|fpga_interfaces|f2h_sdram0_READDATA[54] ;

assign hps_f2h_sdram0_data_readdata[55] = \hps|fpga_interfaces|f2h_sdram0_READDATA[55] ;

assign hps_f2h_sdram0_data_readdata[56] = \hps|fpga_interfaces|f2h_sdram0_READDATA[56] ;

assign hps_f2h_sdram0_data_readdata[57] = \hps|fpga_interfaces|f2h_sdram0_READDATA[57] ;

assign hps_f2h_sdram0_data_readdata[58] = \hps|fpga_interfaces|f2h_sdram0_READDATA[58] ;

assign hps_f2h_sdram0_data_readdata[59] = \hps|fpga_interfaces|f2h_sdram0_READDATA[59] ;

assign hps_f2h_sdram0_data_readdata[60] = \hps|fpga_interfaces|f2h_sdram0_READDATA[60] ;

assign hps_f2h_sdram0_data_readdata[61] = \hps|fpga_interfaces|f2h_sdram0_READDATA[61] ;

assign hps_f2h_sdram0_data_readdata[62] = \hps|fpga_interfaces|f2h_sdram0_READDATA[62] ;

assign hps_f2h_sdram0_data_readdata[63] = \hps|fpga_interfaces|f2h_sdram0_READDATA[63] ;

assign hps_f2h_sdram0_data_readdata[64] = \hps|fpga_interfaces|f2h_sdram0_READDATA[64] ;

assign hps_f2h_sdram0_data_readdata[65] = \hps|fpga_interfaces|f2h_sdram0_READDATA[65] ;

assign hps_f2h_sdram0_data_readdata[66] = \hps|fpga_interfaces|f2h_sdram0_READDATA[66] ;

assign hps_f2h_sdram0_data_readdata[67] = \hps|fpga_interfaces|f2h_sdram0_READDATA[67] ;

assign hps_f2h_sdram0_data_readdata[68] = \hps|fpga_interfaces|f2h_sdram0_READDATA[68] ;

assign hps_f2h_sdram0_data_readdata[69] = \hps|fpga_interfaces|f2h_sdram0_READDATA[69] ;

assign hps_f2h_sdram0_data_readdata[70] = \hps|fpga_interfaces|f2h_sdram0_READDATA[70] ;

assign hps_f2h_sdram0_data_readdata[71] = \hps|fpga_interfaces|f2h_sdram0_READDATA[71] ;

assign hps_f2h_sdram0_data_readdata[72] = \hps|fpga_interfaces|f2h_sdram0_READDATA[72] ;

assign hps_f2h_sdram0_data_readdata[73] = \hps|fpga_interfaces|f2h_sdram0_READDATA[73] ;

assign hps_f2h_sdram0_data_readdata[74] = \hps|fpga_interfaces|f2h_sdram0_READDATA[74] ;

assign hps_f2h_sdram0_data_readdata[75] = \hps|fpga_interfaces|f2h_sdram0_READDATA[75] ;

assign hps_f2h_sdram0_data_readdata[76] = \hps|fpga_interfaces|f2h_sdram0_READDATA[76] ;

assign hps_f2h_sdram0_data_readdata[77] = \hps|fpga_interfaces|f2h_sdram0_READDATA[77] ;

assign hps_f2h_sdram0_data_readdata[78] = \hps|fpga_interfaces|f2h_sdram0_READDATA[78] ;

assign hps_f2h_sdram0_data_readdata[79] = \hps|fpga_interfaces|f2h_sdram0_READDATA[79] ;

assign hps_f2h_sdram0_data_readdata[80] = \hps|fpga_interfaces|f2h_sdram0_READDATA[80] ;

assign hps_f2h_sdram0_data_readdata[81] = \hps|fpga_interfaces|f2h_sdram0_READDATA[81] ;

assign hps_f2h_sdram0_data_readdata[82] = \hps|fpga_interfaces|f2h_sdram0_READDATA[82] ;

assign hps_f2h_sdram0_data_readdata[83] = \hps|fpga_interfaces|f2h_sdram0_READDATA[83] ;

assign hps_f2h_sdram0_data_readdata[84] = \hps|fpga_interfaces|f2h_sdram0_READDATA[84] ;

assign hps_f2h_sdram0_data_readdata[85] = \hps|fpga_interfaces|f2h_sdram0_READDATA[85] ;

assign hps_f2h_sdram0_data_readdata[86] = \hps|fpga_interfaces|f2h_sdram0_READDATA[86] ;

assign hps_f2h_sdram0_data_readdata[87] = \hps|fpga_interfaces|f2h_sdram0_READDATA[87] ;

assign hps_f2h_sdram0_data_readdata[88] = \hps|fpga_interfaces|f2h_sdram0_READDATA[88] ;

assign hps_f2h_sdram0_data_readdata[89] = \hps|fpga_interfaces|f2h_sdram0_READDATA[89] ;

assign hps_f2h_sdram0_data_readdata[90] = \hps|fpga_interfaces|f2h_sdram0_READDATA[90] ;

assign hps_f2h_sdram0_data_readdata[91] = \hps|fpga_interfaces|f2h_sdram0_READDATA[91] ;

assign hps_f2h_sdram0_data_readdata[92] = \hps|fpga_interfaces|f2h_sdram0_READDATA[92] ;

assign hps_f2h_sdram0_data_readdata[93] = \hps|fpga_interfaces|f2h_sdram0_READDATA[93] ;

assign hps_f2h_sdram0_data_readdata[94] = \hps|fpga_interfaces|f2h_sdram0_READDATA[94] ;

assign hps_f2h_sdram0_data_readdata[95] = \hps|fpga_interfaces|f2h_sdram0_READDATA[95] ;

assign hps_f2h_sdram0_data_readdata[96] = \hps|fpga_interfaces|f2h_sdram0_READDATA[96] ;

assign hps_f2h_sdram0_data_readdata[97] = \hps|fpga_interfaces|f2h_sdram0_READDATA[97] ;

assign hps_f2h_sdram0_data_readdata[98] = \hps|fpga_interfaces|f2h_sdram0_READDATA[98] ;

assign hps_f2h_sdram0_data_readdata[99] = \hps|fpga_interfaces|f2h_sdram0_READDATA[99] ;

assign hps_f2h_sdram0_data_readdata[100] = \hps|fpga_interfaces|f2h_sdram0_READDATA[100] ;

assign hps_f2h_sdram0_data_readdata[101] = \hps|fpga_interfaces|f2h_sdram0_READDATA[101] ;

assign hps_f2h_sdram0_data_readdata[102] = \hps|fpga_interfaces|f2h_sdram0_READDATA[102] ;

assign hps_f2h_sdram0_data_readdata[103] = \hps|fpga_interfaces|f2h_sdram0_READDATA[103] ;

assign hps_f2h_sdram0_data_readdata[104] = \hps|fpga_interfaces|f2h_sdram0_READDATA[104] ;

assign hps_f2h_sdram0_data_readdata[105] = \hps|fpga_interfaces|f2h_sdram0_READDATA[105] ;

assign hps_f2h_sdram0_data_readdata[106] = \hps|fpga_interfaces|f2h_sdram0_READDATA[106] ;

assign hps_f2h_sdram0_data_readdata[107] = \hps|fpga_interfaces|f2h_sdram0_READDATA[107] ;

assign hps_f2h_sdram0_data_readdata[108] = \hps|fpga_interfaces|f2h_sdram0_READDATA[108] ;

assign hps_f2h_sdram0_data_readdata[109] = \hps|fpga_interfaces|f2h_sdram0_READDATA[109] ;

assign hps_f2h_sdram0_data_readdata[110] = \hps|fpga_interfaces|f2h_sdram0_READDATA[110] ;

assign hps_f2h_sdram0_data_readdata[111] = \hps|fpga_interfaces|f2h_sdram0_READDATA[111] ;

assign hps_f2h_sdram0_data_readdata[112] = \hps|fpga_interfaces|f2h_sdram0_READDATA[112] ;

assign hps_f2h_sdram0_data_readdata[113] = \hps|fpga_interfaces|f2h_sdram0_READDATA[113] ;

assign hps_f2h_sdram0_data_readdata[114] = \hps|fpga_interfaces|f2h_sdram0_READDATA[114] ;

assign hps_f2h_sdram0_data_readdata[115] = \hps|fpga_interfaces|f2h_sdram0_READDATA[115] ;

assign hps_f2h_sdram0_data_readdata[116] = \hps|fpga_interfaces|f2h_sdram0_READDATA[116] ;

assign hps_f2h_sdram0_data_readdata[117] = \hps|fpga_interfaces|f2h_sdram0_READDATA[117] ;

assign hps_f2h_sdram0_data_readdata[118] = \hps|fpga_interfaces|f2h_sdram0_READDATA[118] ;

assign hps_f2h_sdram0_data_readdata[119] = \hps|fpga_interfaces|f2h_sdram0_READDATA[119] ;

assign hps_f2h_sdram0_data_readdata[120] = \hps|fpga_interfaces|f2h_sdram0_READDATA[120] ;

assign hps_f2h_sdram0_data_readdata[121] = \hps|fpga_interfaces|f2h_sdram0_READDATA[121] ;

assign hps_f2h_sdram0_data_readdata[122] = \hps|fpga_interfaces|f2h_sdram0_READDATA[122] ;

assign hps_f2h_sdram0_data_readdata[123] = \hps|fpga_interfaces|f2h_sdram0_READDATA[123] ;

assign hps_f2h_sdram0_data_readdata[124] = \hps|fpga_interfaces|f2h_sdram0_READDATA[124] ;

assign hps_f2h_sdram0_data_readdata[125] = \hps|fpga_interfaces|f2h_sdram0_READDATA[125] ;

assign hps_f2h_sdram0_data_readdata[126] = \hps|fpga_interfaces|f2h_sdram0_READDATA[126] ;

assign hps_f2h_sdram0_data_readdata[127] = \hps|fpga_interfaces|f2h_sdram0_READDATA[127] ;

assign hps_f2h_sdram0_data_readdata[128] = \hps|fpga_interfaces|f2h_sdram0_READDATA[128] ;

assign hps_f2h_sdram0_data_readdata[129] = \hps|fpga_interfaces|f2h_sdram0_READDATA[129] ;

assign hps_f2h_sdram0_data_readdata[130] = \hps|fpga_interfaces|f2h_sdram0_READDATA[130] ;

assign hps_f2h_sdram0_data_readdata[131] = \hps|fpga_interfaces|f2h_sdram0_READDATA[131] ;

assign hps_f2h_sdram0_data_readdata[132] = \hps|fpga_interfaces|f2h_sdram0_READDATA[132] ;

assign hps_f2h_sdram0_data_readdata[133] = \hps|fpga_interfaces|f2h_sdram0_READDATA[133] ;

assign hps_f2h_sdram0_data_readdata[134] = \hps|fpga_interfaces|f2h_sdram0_READDATA[134] ;

assign hps_f2h_sdram0_data_readdata[135] = \hps|fpga_interfaces|f2h_sdram0_READDATA[135] ;

assign hps_f2h_sdram0_data_readdata[136] = \hps|fpga_interfaces|f2h_sdram0_READDATA[136] ;

assign hps_f2h_sdram0_data_readdata[137] = \hps|fpga_interfaces|f2h_sdram0_READDATA[137] ;

assign hps_f2h_sdram0_data_readdata[138] = \hps|fpga_interfaces|f2h_sdram0_READDATA[138] ;

assign hps_f2h_sdram0_data_readdata[139] = \hps|fpga_interfaces|f2h_sdram0_READDATA[139] ;

assign hps_f2h_sdram0_data_readdata[140] = \hps|fpga_interfaces|f2h_sdram0_READDATA[140] ;

assign hps_f2h_sdram0_data_readdata[141] = \hps|fpga_interfaces|f2h_sdram0_READDATA[141] ;

assign hps_f2h_sdram0_data_readdata[142] = \hps|fpga_interfaces|f2h_sdram0_READDATA[142] ;

assign hps_f2h_sdram0_data_readdata[143] = \hps|fpga_interfaces|f2h_sdram0_READDATA[143] ;

assign hps_f2h_sdram0_data_readdata[144] = \hps|fpga_interfaces|f2h_sdram0_READDATA[144] ;

assign hps_f2h_sdram0_data_readdata[145] = \hps|fpga_interfaces|f2h_sdram0_READDATA[145] ;

assign hps_f2h_sdram0_data_readdata[146] = \hps|fpga_interfaces|f2h_sdram0_READDATA[146] ;

assign hps_f2h_sdram0_data_readdata[147] = \hps|fpga_interfaces|f2h_sdram0_READDATA[147] ;

assign hps_f2h_sdram0_data_readdata[148] = \hps|fpga_interfaces|f2h_sdram0_READDATA[148] ;

assign hps_f2h_sdram0_data_readdata[149] = \hps|fpga_interfaces|f2h_sdram0_READDATA[149] ;

assign hps_f2h_sdram0_data_readdata[150] = \hps|fpga_interfaces|f2h_sdram0_READDATA[150] ;

assign hps_f2h_sdram0_data_readdata[151] = \hps|fpga_interfaces|f2h_sdram0_READDATA[151] ;

assign hps_f2h_sdram0_data_readdata[152] = \hps|fpga_interfaces|f2h_sdram0_READDATA[152] ;

assign hps_f2h_sdram0_data_readdata[153] = \hps|fpga_interfaces|f2h_sdram0_READDATA[153] ;

assign hps_f2h_sdram0_data_readdata[154] = \hps|fpga_interfaces|f2h_sdram0_READDATA[154] ;

assign hps_f2h_sdram0_data_readdata[155] = \hps|fpga_interfaces|f2h_sdram0_READDATA[155] ;

assign hps_f2h_sdram0_data_readdata[156] = \hps|fpga_interfaces|f2h_sdram0_READDATA[156] ;

assign hps_f2h_sdram0_data_readdata[157] = \hps|fpga_interfaces|f2h_sdram0_READDATA[157] ;

assign hps_f2h_sdram0_data_readdata[158] = \hps|fpga_interfaces|f2h_sdram0_READDATA[158] ;

assign hps_f2h_sdram0_data_readdata[159] = \hps|fpga_interfaces|f2h_sdram0_READDATA[159] ;

assign hps_f2h_sdram0_data_readdata[160] = \hps|fpga_interfaces|f2h_sdram0_READDATA[160] ;

assign hps_f2h_sdram0_data_readdata[161] = \hps|fpga_interfaces|f2h_sdram0_READDATA[161] ;

assign hps_f2h_sdram0_data_readdata[162] = \hps|fpga_interfaces|f2h_sdram0_READDATA[162] ;

assign hps_f2h_sdram0_data_readdata[163] = \hps|fpga_interfaces|f2h_sdram0_READDATA[163] ;

assign hps_f2h_sdram0_data_readdata[164] = \hps|fpga_interfaces|f2h_sdram0_READDATA[164] ;

assign hps_f2h_sdram0_data_readdata[165] = \hps|fpga_interfaces|f2h_sdram0_READDATA[165] ;

assign hps_f2h_sdram0_data_readdata[166] = \hps|fpga_interfaces|f2h_sdram0_READDATA[166] ;

assign hps_f2h_sdram0_data_readdata[167] = \hps|fpga_interfaces|f2h_sdram0_READDATA[167] ;

assign hps_f2h_sdram0_data_readdata[168] = \hps|fpga_interfaces|f2h_sdram0_READDATA[168] ;

assign hps_f2h_sdram0_data_readdata[169] = \hps|fpga_interfaces|f2h_sdram0_READDATA[169] ;

assign hps_f2h_sdram0_data_readdata[170] = \hps|fpga_interfaces|f2h_sdram0_READDATA[170] ;

assign hps_f2h_sdram0_data_readdata[171] = \hps|fpga_interfaces|f2h_sdram0_READDATA[171] ;

assign hps_f2h_sdram0_data_readdata[172] = \hps|fpga_interfaces|f2h_sdram0_READDATA[172] ;

assign hps_f2h_sdram0_data_readdata[173] = \hps|fpga_interfaces|f2h_sdram0_READDATA[173] ;

assign hps_f2h_sdram0_data_readdata[174] = \hps|fpga_interfaces|f2h_sdram0_READDATA[174] ;

assign hps_f2h_sdram0_data_readdata[175] = \hps|fpga_interfaces|f2h_sdram0_READDATA[175] ;

assign hps_f2h_sdram0_data_readdata[176] = \hps|fpga_interfaces|f2h_sdram0_READDATA[176] ;

assign hps_f2h_sdram0_data_readdata[177] = \hps|fpga_interfaces|f2h_sdram0_READDATA[177] ;

assign hps_f2h_sdram0_data_readdata[178] = \hps|fpga_interfaces|f2h_sdram0_READDATA[178] ;

assign hps_f2h_sdram0_data_readdata[179] = \hps|fpga_interfaces|f2h_sdram0_READDATA[179] ;

assign hps_f2h_sdram0_data_readdata[180] = \hps|fpga_interfaces|f2h_sdram0_READDATA[180] ;

assign hps_f2h_sdram0_data_readdata[181] = \hps|fpga_interfaces|f2h_sdram0_READDATA[181] ;

assign hps_f2h_sdram0_data_readdata[182] = \hps|fpga_interfaces|f2h_sdram0_READDATA[182] ;

assign hps_f2h_sdram0_data_readdata[183] = \hps|fpga_interfaces|f2h_sdram0_READDATA[183] ;

assign hps_f2h_sdram0_data_readdata[184] = \hps|fpga_interfaces|f2h_sdram0_READDATA[184] ;

assign hps_f2h_sdram0_data_readdata[185] = \hps|fpga_interfaces|f2h_sdram0_READDATA[185] ;

assign hps_f2h_sdram0_data_readdata[186] = \hps|fpga_interfaces|f2h_sdram0_READDATA[186] ;

assign hps_f2h_sdram0_data_readdata[187] = \hps|fpga_interfaces|f2h_sdram0_READDATA[187] ;

assign hps_f2h_sdram0_data_readdata[188] = \hps|fpga_interfaces|f2h_sdram0_READDATA[188] ;

assign hps_f2h_sdram0_data_readdata[189] = \hps|fpga_interfaces|f2h_sdram0_READDATA[189] ;

assign hps_f2h_sdram0_data_readdata[190] = \hps|fpga_interfaces|f2h_sdram0_READDATA[190] ;

assign hps_f2h_sdram0_data_readdata[191] = \hps|fpga_interfaces|f2h_sdram0_READDATA[191] ;

assign hps_f2h_sdram0_data_readdata[192] = \hps|fpga_interfaces|f2h_sdram0_READDATA[192] ;

assign hps_f2h_sdram0_data_readdata[193] = \hps|fpga_interfaces|f2h_sdram0_READDATA[193] ;

assign hps_f2h_sdram0_data_readdata[194] = \hps|fpga_interfaces|f2h_sdram0_READDATA[194] ;

assign hps_f2h_sdram0_data_readdata[195] = \hps|fpga_interfaces|f2h_sdram0_READDATA[195] ;

assign hps_f2h_sdram0_data_readdata[196] = \hps|fpga_interfaces|f2h_sdram0_READDATA[196] ;

assign hps_f2h_sdram0_data_readdata[197] = \hps|fpga_interfaces|f2h_sdram0_READDATA[197] ;

assign hps_f2h_sdram0_data_readdata[198] = \hps|fpga_interfaces|f2h_sdram0_READDATA[198] ;

assign hps_f2h_sdram0_data_readdata[199] = \hps|fpga_interfaces|f2h_sdram0_READDATA[199] ;

assign hps_f2h_sdram0_data_readdata[200] = \hps|fpga_interfaces|f2h_sdram0_READDATA[200] ;

assign hps_f2h_sdram0_data_readdata[201] = \hps|fpga_interfaces|f2h_sdram0_READDATA[201] ;

assign hps_f2h_sdram0_data_readdata[202] = \hps|fpga_interfaces|f2h_sdram0_READDATA[202] ;

assign hps_f2h_sdram0_data_readdata[203] = \hps|fpga_interfaces|f2h_sdram0_READDATA[203] ;

assign hps_f2h_sdram0_data_readdata[204] = \hps|fpga_interfaces|f2h_sdram0_READDATA[204] ;

assign hps_f2h_sdram0_data_readdata[205] = \hps|fpga_interfaces|f2h_sdram0_READDATA[205] ;

assign hps_f2h_sdram0_data_readdata[206] = \hps|fpga_interfaces|f2h_sdram0_READDATA[206] ;

assign hps_f2h_sdram0_data_readdata[207] = \hps|fpga_interfaces|f2h_sdram0_READDATA[207] ;

assign hps_f2h_sdram0_data_readdata[208] = \hps|fpga_interfaces|f2h_sdram0_READDATA[208] ;

assign hps_f2h_sdram0_data_readdata[209] = \hps|fpga_interfaces|f2h_sdram0_READDATA[209] ;

assign hps_f2h_sdram0_data_readdata[210] = \hps|fpga_interfaces|f2h_sdram0_READDATA[210] ;

assign hps_f2h_sdram0_data_readdata[211] = \hps|fpga_interfaces|f2h_sdram0_READDATA[211] ;

assign hps_f2h_sdram0_data_readdata[212] = \hps|fpga_interfaces|f2h_sdram0_READDATA[212] ;

assign hps_f2h_sdram0_data_readdata[213] = \hps|fpga_interfaces|f2h_sdram0_READDATA[213] ;

assign hps_f2h_sdram0_data_readdata[214] = \hps|fpga_interfaces|f2h_sdram0_READDATA[214] ;

assign hps_f2h_sdram0_data_readdata[215] = \hps|fpga_interfaces|f2h_sdram0_READDATA[215] ;

assign hps_f2h_sdram0_data_readdata[216] = \hps|fpga_interfaces|f2h_sdram0_READDATA[216] ;

assign hps_f2h_sdram0_data_readdata[217] = \hps|fpga_interfaces|f2h_sdram0_READDATA[217] ;

assign hps_f2h_sdram0_data_readdata[218] = \hps|fpga_interfaces|f2h_sdram0_READDATA[218] ;

assign hps_f2h_sdram0_data_readdata[219] = \hps|fpga_interfaces|f2h_sdram0_READDATA[219] ;

assign hps_f2h_sdram0_data_readdata[220] = \hps|fpga_interfaces|f2h_sdram0_READDATA[220] ;

assign hps_f2h_sdram0_data_readdata[221] = \hps|fpga_interfaces|f2h_sdram0_READDATA[221] ;

assign hps_f2h_sdram0_data_readdata[222] = \hps|fpga_interfaces|f2h_sdram0_READDATA[222] ;

assign hps_f2h_sdram0_data_readdata[223] = \hps|fpga_interfaces|f2h_sdram0_READDATA[223] ;

assign hps_f2h_sdram0_data_readdata[224] = \hps|fpga_interfaces|f2h_sdram0_READDATA[224] ;

assign hps_f2h_sdram0_data_readdata[225] = \hps|fpga_interfaces|f2h_sdram0_READDATA[225] ;

assign hps_f2h_sdram0_data_readdata[226] = \hps|fpga_interfaces|f2h_sdram0_READDATA[226] ;

assign hps_f2h_sdram0_data_readdata[227] = \hps|fpga_interfaces|f2h_sdram0_READDATA[227] ;

assign hps_f2h_sdram0_data_readdata[228] = \hps|fpga_interfaces|f2h_sdram0_READDATA[228] ;

assign hps_f2h_sdram0_data_readdata[229] = \hps|fpga_interfaces|f2h_sdram0_READDATA[229] ;

assign hps_f2h_sdram0_data_readdata[230] = \hps|fpga_interfaces|f2h_sdram0_READDATA[230] ;

assign hps_f2h_sdram0_data_readdata[231] = \hps|fpga_interfaces|f2h_sdram0_READDATA[231] ;

assign hps_f2h_sdram0_data_readdata[232] = \hps|fpga_interfaces|f2h_sdram0_READDATA[232] ;

assign hps_f2h_sdram0_data_readdata[233] = \hps|fpga_interfaces|f2h_sdram0_READDATA[233] ;

assign hps_f2h_sdram0_data_readdata[234] = \hps|fpga_interfaces|f2h_sdram0_READDATA[234] ;

assign hps_f2h_sdram0_data_readdata[235] = \hps|fpga_interfaces|f2h_sdram0_READDATA[235] ;

assign hps_f2h_sdram0_data_readdata[236] = \hps|fpga_interfaces|f2h_sdram0_READDATA[236] ;

assign hps_f2h_sdram0_data_readdata[237] = \hps|fpga_interfaces|f2h_sdram0_READDATA[237] ;

assign hps_f2h_sdram0_data_readdata[238] = \hps|fpga_interfaces|f2h_sdram0_READDATA[238] ;

assign hps_f2h_sdram0_data_readdata[239] = \hps|fpga_interfaces|f2h_sdram0_READDATA[239] ;

assign hps_f2h_sdram0_data_readdata[240] = \hps|fpga_interfaces|f2h_sdram0_READDATA[240] ;

assign hps_f2h_sdram0_data_readdata[241] = \hps|fpga_interfaces|f2h_sdram0_READDATA[241] ;

assign hps_f2h_sdram0_data_readdata[242] = \hps|fpga_interfaces|f2h_sdram0_READDATA[242] ;

assign hps_f2h_sdram0_data_readdata[243] = \hps|fpga_interfaces|f2h_sdram0_READDATA[243] ;

assign hps_f2h_sdram0_data_readdata[244] = \hps|fpga_interfaces|f2h_sdram0_READDATA[244] ;

assign hps_f2h_sdram0_data_readdata[245] = \hps|fpga_interfaces|f2h_sdram0_READDATA[245] ;

assign hps_f2h_sdram0_data_readdata[246] = \hps|fpga_interfaces|f2h_sdram0_READDATA[246] ;

assign hps_f2h_sdram0_data_readdata[247] = \hps|fpga_interfaces|f2h_sdram0_READDATA[247] ;

assign hps_f2h_sdram0_data_readdata[248] = \hps|fpga_interfaces|f2h_sdram0_READDATA[248] ;

assign hps_f2h_sdram0_data_readdata[249] = \hps|fpga_interfaces|f2h_sdram0_READDATA[249] ;

assign hps_f2h_sdram0_data_readdata[250] = \hps|fpga_interfaces|f2h_sdram0_READDATA[250] ;

assign hps_f2h_sdram0_data_readdata[251] = \hps|fpga_interfaces|f2h_sdram0_READDATA[251] ;

assign hps_f2h_sdram0_data_readdata[252] = \hps|fpga_interfaces|f2h_sdram0_READDATA[252] ;

assign hps_f2h_sdram0_data_readdata[253] = \hps|fpga_interfaces|f2h_sdram0_READDATA[253] ;

assign hps_f2h_sdram0_data_readdata[254] = \hps|fpga_interfaces|f2h_sdram0_READDATA[254] ;

assign hps_f2h_sdram0_data_readdata[255] = \hps|fpga_interfaces|f2h_sdram0_READDATA[255] ;

assign hps_f2h_sdram0_data_readdatavalid = \hps|fpga_interfaces|f2h_sdram0_READDATAVALID[0] ;

assign hps_h2f_cold_reset_reset_n = \hps|fpga_interfaces|h2f_cold_rst_n[0] ;

assign hps_h2f_warm_reset_handshake_h2f_pending_rst_req_n = \hps|fpga_interfaces|h2f_pending_rst_req_n[0] ;

assign hps_hps_io_hps_io_emac1_inst_TX_CLK = \hps|hps_io|border|emac1_inst~O_EMAC_CLK_TX ;

assign hps_hps_io_hps_io_emac1_inst_TXD0 = \hps|hps_io|border|emac1_inst~emac_phy_txd ;

assign hps_hps_io_hps_io_emac1_inst_TXD1 = \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD1 ;

assign hps_hps_io_hps_io_emac1_inst_TXD2 = \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD2 ;

assign hps_hps_io_hps_io_emac1_inst_TXD3 = \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TXD3 ;

assign hps_hps_io_hps_io_emac1_inst_MDC = \hps|hps_io|border|emac1_inst~O_EMAC_GMII_MDC ;

assign hps_hps_io_hps_io_emac1_inst_TX_CTL = \hps|hps_io|border|emac1_inst~O_EMAC_PHY_TX_OE ;

assign hps_hps_io_hps_io_sdio_inst_CLK = \hps|hps_io|border|sdio_inst~sdmmc_cclk ;

assign hps_hps_io_hps_io_uart0_inst_TX = \hps|hps_io|border|uart0_inst~uart_txd ;

assign leds_out_export[0] = \leds|data_out[0]~q ;

assign leds_out_export[1] = \leds|data_out[1]~q ;

assign leds_out_export[2] = \leds|data_out[2]~q ;

assign leds_out_export[3] = \leds|data_out[3]~q ;

assign leds_out_export[4] = \leds|data_out[4]~q ;

assign leds_out_export[5] = \leds|data_out[5]~q ;

assign leds_out_export[6] = \leds|data_out[6]~q ;

assign leds_out_export[7] = \leds|data_out[7]~q ;

assign leds_out_export[8] = \leds|data_out[8]~q ;

assign leds_out_export[9] = \leds|data_out[9]~q ;

assign memory_mem_a[0] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[0] ;

assign memory_mem_a[1] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[1] ;

assign memory_mem_a[2] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[2] ;

assign memory_mem_a[3] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[3] ;

assign memory_mem_a[4] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[4] ;

assign memory_mem_a[5] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[5] ;

assign memory_mem_a[6] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[6] ;

assign memory_mem_a[7] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[7] ;

assign memory_mem_a[8] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[8] ;

assign memory_mem_a[9] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[9] ;

assign memory_mem_a[10] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[10] ;

assign memory_mem_a[11] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[11] ;

assign memory_mem_a[12] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[12] ;

assign memory_mem_a[13] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[13] ;

assign memory_mem_a[14] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|uaddress_pad|dataout[14] ;

assign memory_mem_ba[0] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[0] ;

assign memory_mem_ba[1] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[1] ;

assign memory_mem_ba[2] = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ubank_pad|dataout[2] ;

assign memory_mem_cke = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[1] ;

assign memory_mem_cs_n = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[0] ;

assign memory_mem_ras_n = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[3] ;

assign memory_mem_cas_n = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[4] ;

assign memory_mem_we_n = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[5] ;

assign memory_mem_reset_n = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ureset_n_pad|dataout[0] ;

assign memory_mem_odt = \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|uaddr_cmd_pads|ucmd_pad|dataout[2] ;

cyclonev_io_obuf \hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output (
	.i(\hps|hps_io|border|intermediate[0] ),
	.oe(\hps|hps_io|border|intermediate[1] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_hps_io_hps_io_emac1_inst_MDIO),
	.obar());
defparam \hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .bus_hold = "false";
defparam \hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .open_drain_output = "false";
defparam \hps|hps_io|border|hps_io_emac1_inst_MDIO[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output (
	.i(\hps|hps_io|border|intermediate[2] ),
	.oe(\hps|hps_io|border|intermediate[3] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_hps_io_hps_io_sdio_inst_CMD),
	.obar());
defparam \hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .bus_hold = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .open_drain_output = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_CMD[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_io_sdio_inst_D0[0]~output (
	.i(\hps|hps_io|border|intermediate[4] ),
	.oe(\hps|hps_io|border|intermediate[5] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_hps_io_hps_io_sdio_inst_D0),
	.obar());
defparam \hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .bus_hold = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .open_drain_output = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D0[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_io_sdio_inst_D1[0]~output (
	.i(\hps|hps_io|border|intermediate[6] ),
	.oe(\hps|hps_io|border|intermediate[7] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_hps_io_hps_io_sdio_inst_D1),
	.obar());
defparam \hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .bus_hold = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .open_drain_output = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D1[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_io_sdio_inst_D2[0]~output (
	.i(\hps|hps_io|border|intermediate[8] ),
	.oe(\hps|hps_io|border|intermediate[9] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_hps_io_hps_io_sdio_inst_D2),
	.obar());
defparam \hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .bus_hold = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .open_drain_output = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D2[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_io_sdio_inst_D3[0]~output (
	.i(\hps|hps_io|border|intermediate[10] ),
	.oe(\hps|hps_io|border|intermediate[11] ),
	.dynamicterminationcontrol(gnd),
	.seriesterminationcontrol(16'b0000000000000000),
	.parallelterminationcontrol(16'b0000000000000000),
	.o(hps_hps_io_hps_io_sdio_inst_D3),
	.obar());
defparam \hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .bus_hold = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .open_drain_output = "false";
defparam \hps|hps_io|border|hps_io_sdio_inst_D3[0]~output .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[0]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[1]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[2]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[3]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[4]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[5]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[6]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[7]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[8]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[9]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[10]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[11]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[12]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[13]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[14]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[15]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[16]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[17]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[18]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[19]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[20]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[21]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[22]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[23]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[24]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[0].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[25]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[1].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[26]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[2].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[27]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[3].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[28]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[4].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[29]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[5].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[30]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[6].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_data_out ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].delayed_oe_1 ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|delayed_oct ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dq[31]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|pad_gen[7].data_out .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[0]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[1]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[2]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs[3]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[0]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[1]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[2]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

cyclonev_io_obuf \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 (
	.i(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|os_bar ),
	.oe(!\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_oe_bar ),
	.dynamicterminationcontrol(\hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|diff_dtc_bar ),
	.seriesterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|seriesterminationcontrol[0] }),
	.parallelterminationcontrol({\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[15] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[14] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[13] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[12] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[11] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[10] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[9] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[8] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[7] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[6] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[5] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[4] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[3] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[2] ,\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[1] ,
\hps|hps_io|border|hps_sdram_inst|oct|parallelterminationcontrol[0] }),
	.o(memory_mem_dqs_n[3]),
	.obar());
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .bus_hold = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .open_drain_output = "false";
defparam \hps|hps_io|border|hps_sdram_inst|p0|umemphy|uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|obuf_os_bar_0 .shift_series_termination_control = "false";

endmodule

module terminal_qsys_terminal_qsys_base_address_ddr (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	data_out_24,
	data_out_25,
	data_out_26,
	data_out_27,
	data_out_28,
	data_out_29,
	data_out_30,
	data_out_31,
	wait_latency_counter_1,
	wait_latency_counter_0,
	writedata,
	reset_n,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	readdata_18,
	readdata_19,
	readdata_20,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_16;
output 	data_out_17;
output 	data_out_18;
output 	data_out_19;
output 	data_out_20;
output 	data_out_21;
output 	data_out_22;
output 	data_out_23;
output 	data_out_24;
output 	data_out_25;
output 	data_out_26;
output 	data_out_27;
output 	data_out_28;
output 	data_out_29;
output 	data_out_30;
output 	data_out_31;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	[31:0] writedata;
input 	reset_n;
input 	m0_write;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
output 	readdata_18;
output 	readdata_19;
output 	readdata_20;
output 	readdata_21;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(writedata[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(writedata[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \data_out[18] (
	.clk(clk),
	.d(writedata[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_18),
	.prn(vcc));
defparam \data_out[18] .is_wysiwyg = "true";
defparam \data_out[18] .power_up = "low";

dffeas \data_out[19] (
	.clk(clk),
	.d(writedata[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_19),
	.prn(vcc));
defparam \data_out[19] .is_wysiwyg = "true";
defparam \data_out[19] .power_up = "low";

dffeas \data_out[20] (
	.clk(clk),
	.d(writedata[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_20),
	.prn(vcc));
defparam \data_out[20] .is_wysiwyg = "true";
defparam \data_out[20] .power_up = "low";

dffeas \data_out[21] (
	.clk(clk),
	.d(writedata[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_21),
	.prn(vcc));
defparam \data_out[21] .is_wysiwyg = "true";
defparam \data_out[21] .power_up = "low";

dffeas \data_out[22] (
	.clk(clk),
	.d(writedata[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_22),
	.prn(vcc));
defparam \data_out[22] .is_wysiwyg = "true";
defparam \data_out[22] .power_up = "low";

dffeas \data_out[23] (
	.clk(clk),
	.d(writedata[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_23),
	.prn(vcc));
defparam \data_out[23] .is_wysiwyg = "true";
defparam \data_out[23] .power_up = "low";

dffeas \data_out[24] (
	.clk(clk),
	.d(writedata[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_24),
	.prn(vcc));
defparam \data_out[24] .is_wysiwyg = "true";
defparam \data_out[24] .power_up = "low";

dffeas \data_out[25] (
	.clk(clk),
	.d(writedata[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_25),
	.prn(vcc));
defparam \data_out[25] .is_wysiwyg = "true";
defparam \data_out[25] .power_up = "low";

dffeas \data_out[26] (
	.clk(clk),
	.d(writedata[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_26),
	.prn(vcc));
defparam \data_out[26] .is_wysiwyg = "true";
defparam \data_out[26] .power_up = "low";

dffeas \data_out[27] (
	.clk(clk),
	.d(writedata[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_27),
	.prn(vcc));
defparam \data_out[27] .is_wysiwyg = "true";
defparam \data_out[27] .power_up = "low";

dffeas \data_out[28] (
	.clk(clk),
	.d(writedata[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_28),
	.prn(vcc));
defparam \data_out[28] .is_wysiwyg = "true";
defparam \data_out[28] .power_up = "low";

dffeas \data_out[29] (
	.clk(clk),
	.d(writedata[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_29),
	.prn(vcc));
defparam \data_out[29] .is_wysiwyg = "true";
defparam \data_out[29] .power_up = "low";

dffeas \data_out[30] (
	.clk(clk),
	.d(writedata[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_30),
	.prn(vcc));
defparam \data_out[30] .is_wysiwyg = "true";
defparam \data_out[30] .power_up = "low";

dffeas \data_out[31] (
	.clk(clk),
	.d(writedata[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_31),
	.prn(vcc));
defparam \data_out[31] .is_wysiwyg = "true";
defparam \data_out[31] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'h4040404040404040;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'h4040404040404040;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'h4040404040404040;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'h4040404040404040;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'h4040404040404040;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'h4040404040404040;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'h4040404040404040;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'h4040404040404040;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \readdata[8] (
	.dataa(!data_out_8),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[8] .extended_lut = "off";
defparam \readdata[8] .lut_mask = 64'h4040404040404040;
defparam \readdata[8] .shared_arith = "off";

cyclonev_lcell_comb \readdata[9] (
	.dataa(!data_out_9),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[9] .extended_lut = "off";
defparam \readdata[9] .lut_mask = 64'h4040404040404040;
defparam \readdata[9] .shared_arith = "off";

cyclonev_lcell_comb \readdata[10] (
	.dataa(!data_out_10),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[10] .extended_lut = "off";
defparam \readdata[10] .lut_mask = 64'h4040404040404040;
defparam \readdata[10] .shared_arith = "off";

cyclonev_lcell_comb \readdata[11] (
	.dataa(!data_out_11),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[11] .extended_lut = "off";
defparam \readdata[11] .lut_mask = 64'h4040404040404040;
defparam \readdata[11] .shared_arith = "off";

cyclonev_lcell_comb \readdata[12] (
	.dataa(!data_out_12),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[12] .extended_lut = "off";
defparam \readdata[12] .lut_mask = 64'h4040404040404040;
defparam \readdata[12] .shared_arith = "off";

cyclonev_lcell_comb \readdata[13] (
	.dataa(!data_out_13),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[13] .extended_lut = "off";
defparam \readdata[13] .lut_mask = 64'h4040404040404040;
defparam \readdata[13] .shared_arith = "off";

cyclonev_lcell_comb \readdata[14] (
	.dataa(!data_out_14),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[14] .extended_lut = "off";
defparam \readdata[14] .lut_mask = 64'h4040404040404040;
defparam \readdata[14] .shared_arith = "off";

cyclonev_lcell_comb \readdata[15] (
	.dataa(!data_out_15),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[15] .extended_lut = "off";
defparam \readdata[15] .lut_mask = 64'h4040404040404040;
defparam \readdata[15] .shared_arith = "off";

cyclonev_lcell_comb \readdata[16] (
	.dataa(!data_out_16),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[16] .extended_lut = "off";
defparam \readdata[16] .lut_mask = 64'h4040404040404040;
defparam \readdata[16] .shared_arith = "off";

cyclonev_lcell_comb \readdata[17] (
	.dataa(!data_out_17),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[17] .extended_lut = "off";
defparam \readdata[17] .lut_mask = 64'h4040404040404040;
defparam \readdata[17] .shared_arith = "off";

cyclonev_lcell_comb \readdata[18] (
	.dataa(!data_out_18),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[18] .extended_lut = "off";
defparam \readdata[18] .lut_mask = 64'h4040404040404040;
defparam \readdata[18] .shared_arith = "off";

cyclonev_lcell_comb \readdata[19] (
	.dataa(!data_out_19),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[19] .extended_lut = "off";
defparam \readdata[19] .lut_mask = 64'h4040404040404040;
defparam \readdata[19] .shared_arith = "off";

cyclonev_lcell_comb \readdata[20] (
	.dataa(!data_out_20),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[20] .extended_lut = "off";
defparam \readdata[20] .lut_mask = 64'h4040404040404040;
defparam \readdata[20] .shared_arith = "off";

cyclonev_lcell_comb \readdata[21] (
	.dataa(!data_out_21),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[21] .extended_lut = "off";
defparam \readdata[21] .lut_mask = 64'h4040404040404040;
defparam \readdata[21] .shared_arith = "off";

cyclonev_lcell_comb \readdata[22] (
	.dataa(!data_out_22),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[22] .extended_lut = "off";
defparam \readdata[22] .lut_mask = 64'h4040404040404040;
defparam \readdata[22] .shared_arith = "off";

cyclonev_lcell_comb \readdata[23] (
	.dataa(!data_out_23),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[23] .extended_lut = "off";
defparam \readdata[23] .lut_mask = 64'h4040404040404040;
defparam \readdata[23] .shared_arith = "off";

cyclonev_lcell_comb \readdata[24] (
	.dataa(!data_out_24),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[24] .extended_lut = "off";
defparam \readdata[24] .lut_mask = 64'h4040404040404040;
defparam \readdata[24] .shared_arith = "off";

cyclonev_lcell_comb \readdata[25] (
	.dataa(!data_out_25),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[25] .extended_lut = "off";
defparam \readdata[25] .lut_mask = 64'h4040404040404040;
defparam \readdata[25] .shared_arith = "off";

cyclonev_lcell_comb \readdata[26] (
	.dataa(!data_out_26),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[26] .extended_lut = "off";
defparam \readdata[26] .lut_mask = 64'h4040404040404040;
defparam \readdata[26] .shared_arith = "off";

cyclonev_lcell_comb \readdata[27] (
	.dataa(!data_out_27),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[27] .extended_lut = "off";
defparam \readdata[27] .lut_mask = 64'h4040404040404040;
defparam \readdata[27] .shared_arith = "off";

cyclonev_lcell_comb \readdata[28] (
	.dataa(!data_out_28),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[28] .extended_lut = "off";
defparam \readdata[28] .lut_mask = 64'h4040404040404040;
defparam \readdata[28] .shared_arith = "off";

cyclonev_lcell_comb \readdata[29] (
	.dataa(!data_out_29),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[29] .extended_lut = "off";
defparam \readdata[29] .lut_mask = 64'h4040404040404040;
defparam \readdata[29] .shared_arith = "off";

cyclonev_lcell_comb \readdata[30] (
	.dataa(!data_out_30),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[30] .extended_lut = "off";
defparam \readdata[30] .lut_mask = 64'h4040404040404040;
defparam \readdata[30] .shared_arith = "off";

cyclonev_lcell_comb \readdata[31] (
	.dataa(!data_out_31),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[31] .extended_lut = "off";
defparam \readdata[31] .lut_mask = 64'h4040404040404040;
defparam \readdata[31] .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0800000008000000;
defparam \always0~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_base_address_ddr_1 (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	data_out_24,
	data_out_25,
	data_out_26,
	data_out_27,
	data_out_28,
	data_out_29,
	data_out_30,
	data_out_31,
	wait_latency_counter_1,
	wait_latency_counter_0,
	writedata,
	reset_n,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	readdata_18,
	readdata_19,
	readdata_20,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_16;
output 	data_out_17;
output 	data_out_18;
output 	data_out_19;
output 	data_out_20;
output 	data_out_21;
output 	data_out_22;
output 	data_out_23;
output 	data_out_24;
output 	data_out_25;
output 	data_out_26;
output 	data_out_27;
output 	data_out_28;
output 	data_out_29;
output 	data_out_30;
output 	data_out_31;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	[31:0] writedata;
input 	reset_n;
input 	m0_write;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
output 	readdata_18;
output 	readdata_19;
output 	readdata_20;
output 	readdata_21;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(writedata[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(writedata[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \data_out[18] (
	.clk(clk),
	.d(writedata[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_18),
	.prn(vcc));
defparam \data_out[18] .is_wysiwyg = "true";
defparam \data_out[18] .power_up = "low";

dffeas \data_out[19] (
	.clk(clk),
	.d(writedata[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_19),
	.prn(vcc));
defparam \data_out[19] .is_wysiwyg = "true";
defparam \data_out[19] .power_up = "low";

dffeas \data_out[20] (
	.clk(clk),
	.d(writedata[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_20),
	.prn(vcc));
defparam \data_out[20] .is_wysiwyg = "true";
defparam \data_out[20] .power_up = "low";

dffeas \data_out[21] (
	.clk(clk),
	.d(writedata[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_21),
	.prn(vcc));
defparam \data_out[21] .is_wysiwyg = "true";
defparam \data_out[21] .power_up = "low";

dffeas \data_out[22] (
	.clk(clk),
	.d(writedata[22]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_22),
	.prn(vcc));
defparam \data_out[22] .is_wysiwyg = "true";
defparam \data_out[22] .power_up = "low";

dffeas \data_out[23] (
	.clk(clk),
	.d(writedata[23]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_23),
	.prn(vcc));
defparam \data_out[23] .is_wysiwyg = "true";
defparam \data_out[23] .power_up = "low";

dffeas \data_out[24] (
	.clk(clk),
	.d(writedata[24]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_24),
	.prn(vcc));
defparam \data_out[24] .is_wysiwyg = "true";
defparam \data_out[24] .power_up = "low";

dffeas \data_out[25] (
	.clk(clk),
	.d(writedata[25]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_25),
	.prn(vcc));
defparam \data_out[25] .is_wysiwyg = "true";
defparam \data_out[25] .power_up = "low";

dffeas \data_out[26] (
	.clk(clk),
	.d(writedata[26]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_26),
	.prn(vcc));
defparam \data_out[26] .is_wysiwyg = "true";
defparam \data_out[26] .power_up = "low";

dffeas \data_out[27] (
	.clk(clk),
	.d(writedata[27]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_27),
	.prn(vcc));
defparam \data_out[27] .is_wysiwyg = "true";
defparam \data_out[27] .power_up = "low";

dffeas \data_out[28] (
	.clk(clk),
	.d(writedata[28]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_28),
	.prn(vcc));
defparam \data_out[28] .is_wysiwyg = "true";
defparam \data_out[28] .power_up = "low";

dffeas \data_out[29] (
	.clk(clk),
	.d(writedata[29]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_29),
	.prn(vcc));
defparam \data_out[29] .is_wysiwyg = "true";
defparam \data_out[29] .power_up = "low";

dffeas \data_out[30] (
	.clk(clk),
	.d(writedata[30]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_30),
	.prn(vcc));
defparam \data_out[30] .is_wysiwyg = "true";
defparam \data_out[30] .power_up = "low";

dffeas \data_out[31] (
	.clk(clk),
	.d(writedata[31]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_31),
	.prn(vcc));
defparam \data_out[31] .is_wysiwyg = "true";
defparam \data_out[31] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'h4040404040404040;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'h4040404040404040;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'h4040404040404040;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'h4040404040404040;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'h4040404040404040;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'h4040404040404040;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'h4040404040404040;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'h4040404040404040;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \readdata[8] (
	.dataa(!data_out_8),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[8] .extended_lut = "off";
defparam \readdata[8] .lut_mask = 64'h4040404040404040;
defparam \readdata[8] .shared_arith = "off";

cyclonev_lcell_comb \readdata[9] (
	.dataa(!data_out_9),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[9] .extended_lut = "off";
defparam \readdata[9] .lut_mask = 64'h4040404040404040;
defparam \readdata[9] .shared_arith = "off";

cyclonev_lcell_comb \readdata[10] (
	.dataa(!data_out_10),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[10] .extended_lut = "off";
defparam \readdata[10] .lut_mask = 64'h4040404040404040;
defparam \readdata[10] .shared_arith = "off";

cyclonev_lcell_comb \readdata[11] (
	.dataa(!data_out_11),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[11] .extended_lut = "off";
defparam \readdata[11] .lut_mask = 64'h4040404040404040;
defparam \readdata[11] .shared_arith = "off";

cyclonev_lcell_comb \readdata[12] (
	.dataa(!data_out_12),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[12] .extended_lut = "off";
defparam \readdata[12] .lut_mask = 64'h4040404040404040;
defparam \readdata[12] .shared_arith = "off";

cyclonev_lcell_comb \readdata[13] (
	.dataa(!data_out_13),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[13] .extended_lut = "off";
defparam \readdata[13] .lut_mask = 64'h4040404040404040;
defparam \readdata[13] .shared_arith = "off";

cyclonev_lcell_comb \readdata[14] (
	.dataa(!data_out_14),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[14] .extended_lut = "off";
defparam \readdata[14] .lut_mask = 64'h4040404040404040;
defparam \readdata[14] .shared_arith = "off";

cyclonev_lcell_comb \readdata[15] (
	.dataa(!data_out_15),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[15] .extended_lut = "off";
defparam \readdata[15] .lut_mask = 64'h4040404040404040;
defparam \readdata[15] .shared_arith = "off";

cyclonev_lcell_comb \readdata[16] (
	.dataa(!data_out_16),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[16] .extended_lut = "off";
defparam \readdata[16] .lut_mask = 64'h4040404040404040;
defparam \readdata[16] .shared_arith = "off";

cyclonev_lcell_comb \readdata[17] (
	.dataa(!data_out_17),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[17] .extended_lut = "off";
defparam \readdata[17] .lut_mask = 64'h4040404040404040;
defparam \readdata[17] .shared_arith = "off";

cyclonev_lcell_comb \readdata[18] (
	.dataa(!data_out_18),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[18] .extended_lut = "off";
defparam \readdata[18] .lut_mask = 64'h4040404040404040;
defparam \readdata[18] .shared_arith = "off";

cyclonev_lcell_comb \readdata[19] (
	.dataa(!data_out_19),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[19] .extended_lut = "off";
defparam \readdata[19] .lut_mask = 64'h4040404040404040;
defparam \readdata[19] .shared_arith = "off";

cyclonev_lcell_comb \readdata[20] (
	.dataa(!data_out_20),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[20] .extended_lut = "off";
defparam \readdata[20] .lut_mask = 64'h4040404040404040;
defparam \readdata[20] .shared_arith = "off";

cyclonev_lcell_comb \readdata[21] (
	.dataa(!data_out_21),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[21] .extended_lut = "off";
defparam \readdata[21] .lut_mask = 64'h4040404040404040;
defparam \readdata[21] .shared_arith = "off";

cyclonev_lcell_comb \readdata[22] (
	.dataa(!data_out_22),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[22] .extended_lut = "off";
defparam \readdata[22] .lut_mask = 64'h4040404040404040;
defparam \readdata[22] .shared_arith = "off";

cyclonev_lcell_comb \readdata[23] (
	.dataa(!data_out_23),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[23] .extended_lut = "off";
defparam \readdata[23] .lut_mask = 64'h4040404040404040;
defparam \readdata[23] .shared_arith = "off";

cyclonev_lcell_comb \readdata[24] (
	.dataa(!data_out_24),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[24] .extended_lut = "off";
defparam \readdata[24] .lut_mask = 64'h4040404040404040;
defparam \readdata[24] .shared_arith = "off";

cyclonev_lcell_comb \readdata[25] (
	.dataa(!data_out_25),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[25] .extended_lut = "off";
defparam \readdata[25] .lut_mask = 64'h4040404040404040;
defparam \readdata[25] .shared_arith = "off";

cyclonev_lcell_comb \readdata[26] (
	.dataa(!data_out_26),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[26] .extended_lut = "off";
defparam \readdata[26] .lut_mask = 64'h4040404040404040;
defparam \readdata[26] .shared_arith = "off";

cyclonev_lcell_comb \readdata[27] (
	.dataa(!data_out_27),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[27] .extended_lut = "off";
defparam \readdata[27] .lut_mask = 64'h4040404040404040;
defparam \readdata[27] .shared_arith = "off";

cyclonev_lcell_comb \readdata[28] (
	.dataa(!data_out_28),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[28] .extended_lut = "off";
defparam \readdata[28] .lut_mask = 64'h4040404040404040;
defparam \readdata[28] .shared_arith = "off";

cyclonev_lcell_comb \readdata[29] (
	.dataa(!data_out_29),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[29] .extended_lut = "off";
defparam \readdata[29] .lut_mask = 64'h4040404040404040;
defparam \readdata[29] .shared_arith = "off";

cyclonev_lcell_comb \readdata[30] (
	.dataa(!data_out_30),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[30] .extended_lut = "off";
defparam \readdata[30] .lut_mask = 64'h4040404040404040;
defparam \readdata[30] .shared_arith = "off";

cyclonev_lcell_comb \readdata[31] (
	.dataa(!data_out_31),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[31] .extended_lut = "off";
defparam \readdata[31] .lut_mask = 64'h4040404040404040;
defparam \readdata[31] .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0800000008000000;
defparam \always0~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_hps (
	h2f_cold_rst_n_0,
	h2f_pending_rst_req_n_0,
	h2f_rst_n_0,
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARADDR_15,
	h2f_lw_ARADDR_16,
	h2f_lw_ARADDR_17,
	h2f_lw_ARADDR_18,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWADDR_15,
	h2f_lw_AWADDR_16,
	h2f_lw_AWADDR_17,
	h2f_lw_AWADDR_18,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	intermediate_1,
	f2h_sdram0_READDATAVALID_0,
	f2h_sdram0_READDATA_0,
	f2h_sdram0_READDATA_1,
	f2h_sdram0_READDATA_2,
	f2h_sdram0_READDATA_3,
	f2h_sdram0_READDATA_4,
	f2h_sdram0_READDATA_5,
	f2h_sdram0_READDATA_6,
	f2h_sdram0_READDATA_7,
	f2h_sdram0_READDATA_8,
	f2h_sdram0_READDATA_9,
	f2h_sdram0_READDATA_10,
	f2h_sdram0_READDATA_11,
	f2h_sdram0_READDATA_12,
	f2h_sdram0_READDATA_13,
	f2h_sdram0_READDATA_14,
	f2h_sdram0_READDATA_15,
	f2h_sdram0_READDATA_16,
	f2h_sdram0_READDATA_17,
	f2h_sdram0_READDATA_18,
	f2h_sdram0_READDATA_19,
	f2h_sdram0_READDATA_20,
	f2h_sdram0_READDATA_21,
	f2h_sdram0_READDATA_22,
	f2h_sdram0_READDATA_23,
	f2h_sdram0_READDATA_24,
	f2h_sdram0_READDATA_25,
	f2h_sdram0_READDATA_26,
	f2h_sdram0_READDATA_27,
	f2h_sdram0_READDATA_28,
	f2h_sdram0_READDATA_29,
	f2h_sdram0_READDATA_30,
	f2h_sdram0_READDATA_31,
	f2h_sdram0_READDATA_32,
	f2h_sdram0_READDATA_33,
	f2h_sdram0_READDATA_34,
	f2h_sdram0_READDATA_35,
	f2h_sdram0_READDATA_36,
	f2h_sdram0_READDATA_37,
	f2h_sdram0_READDATA_38,
	f2h_sdram0_READDATA_39,
	f2h_sdram0_READDATA_40,
	f2h_sdram0_READDATA_41,
	f2h_sdram0_READDATA_42,
	f2h_sdram0_READDATA_43,
	f2h_sdram0_READDATA_44,
	f2h_sdram0_READDATA_45,
	f2h_sdram0_READDATA_46,
	f2h_sdram0_READDATA_47,
	f2h_sdram0_READDATA_48,
	f2h_sdram0_READDATA_49,
	f2h_sdram0_READDATA_50,
	f2h_sdram0_READDATA_51,
	f2h_sdram0_READDATA_52,
	f2h_sdram0_READDATA_53,
	f2h_sdram0_READDATA_54,
	f2h_sdram0_READDATA_55,
	f2h_sdram0_READDATA_56,
	f2h_sdram0_READDATA_57,
	f2h_sdram0_READDATA_58,
	f2h_sdram0_READDATA_59,
	f2h_sdram0_READDATA_60,
	f2h_sdram0_READDATA_61,
	f2h_sdram0_READDATA_62,
	f2h_sdram0_READDATA_63,
	f2h_sdram0_READDATA_64,
	f2h_sdram0_READDATA_65,
	f2h_sdram0_READDATA_66,
	f2h_sdram0_READDATA_67,
	f2h_sdram0_READDATA_68,
	f2h_sdram0_READDATA_69,
	f2h_sdram0_READDATA_70,
	f2h_sdram0_READDATA_71,
	f2h_sdram0_READDATA_72,
	f2h_sdram0_READDATA_73,
	f2h_sdram0_READDATA_74,
	f2h_sdram0_READDATA_75,
	f2h_sdram0_READDATA_76,
	f2h_sdram0_READDATA_77,
	f2h_sdram0_READDATA_78,
	f2h_sdram0_READDATA_79,
	f2h_sdram0_READDATA_80,
	f2h_sdram0_READDATA_81,
	f2h_sdram0_READDATA_82,
	f2h_sdram0_READDATA_83,
	f2h_sdram0_READDATA_84,
	f2h_sdram0_READDATA_85,
	f2h_sdram0_READDATA_86,
	f2h_sdram0_READDATA_87,
	f2h_sdram0_READDATA_88,
	f2h_sdram0_READDATA_89,
	f2h_sdram0_READDATA_90,
	f2h_sdram0_READDATA_91,
	f2h_sdram0_READDATA_92,
	f2h_sdram0_READDATA_93,
	f2h_sdram0_READDATA_94,
	f2h_sdram0_READDATA_95,
	f2h_sdram0_READDATA_96,
	f2h_sdram0_READDATA_97,
	f2h_sdram0_READDATA_98,
	f2h_sdram0_READDATA_99,
	f2h_sdram0_READDATA_100,
	f2h_sdram0_READDATA_101,
	f2h_sdram0_READDATA_102,
	f2h_sdram0_READDATA_103,
	f2h_sdram0_READDATA_104,
	f2h_sdram0_READDATA_105,
	f2h_sdram0_READDATA_106,
	f2h_sdram0_READDATA_107,
	f2h_sdram0_READDATA_108,
	f2h_sdram0_READDATA_109,
	f2h_sdram0_READDATA_110,
	f2h_sdram0_READDATA_111,
	f2h_sdram0_READDATA_112,
	f2h_sdram0_READDATA_113,
	f2h_sdram0_READDATA_114,
	f2h_sdram0_READDATA_115,
	f2h_sdram0_READDATA_116,
	f2h_sdram0_READDATA_117,
	f2h_sdram0_READDATA_118,
	f2h_sdram0_READDATA_119,
	f2h_sdram0_READDATA_120,
	f2h_sdram0_READDATA_121,
	f2h_sdram0_READDATA_122,
	f2h_sdram0_READDATA_123,
	f2h_sdram0_READDATA_124,
	f2h_sdram0_READDATA_125,
	f2h_sdram0_READDATA_126,
	f2h_sdram0_READDATA_127,
	f2h_sdram0_READDATA_128,
	f2h_sdram0_READDATA_129,
	f2h_sdram0_READDATA_130,
	f2h_sdram0_READDATA_131,
	f2h_sdram0_READDATA_132,
	f2h_sdram0_READDATA_133,
	f2h_sdram0_READDATA_134,
	f2h_sdram0_READDATA_135,
	f2h_sdram0_READDATA_136,
	f2h_sdram0_READDATA_137,
	f2h_sdram0_READDATA_138,
	f2h_sdram0_READDATA_139,
	f2h_sdram0_READDATA_140,
	f2h_sdram0_READDATA_141,
	f2h_sdram0_READDATA_142,
	f2h_sdram0_READDATA_143,
	f2h_sdram0_READDATA_144,
	f2h_sdram0_READDATA_145,
	f2h_sdram0_READDATA_146,
	f2h_sdram0_READDATA_147,
	f2h_sdram0_READDATA_148,
	f2h_sdram0_READDATA_149,
	f2h_sdram0_READDATA_150,
	f2h_sdram0_READDATA_151,
	f2h_sdram0_READDATA_152,
	f2h_sdram0_READDATA_153,
	f2h_sdram0_READDATA_154,
	f2h_sdram0_READDATA_155,
	f2h_sdram0_READDATA_156,
	f2h_sdram0_READDATA_157,
	f2h_sdram0_READDATA_158,
	f2h_sdram0_READDATA_159,
	f2h_sdram0_READDATA_160,
	f2h_sdram0_READDATA_161,
	f2h_sdram0_READDATA_162,
	f2h_sdram0_READDATA_163,
	f2h_sdram0_READDATA_164,
	f2h_sdram0_READDATA_165,
	f2h_sdram0_READDATA_166,
	f2h_sdram0_READDATA_167,
	f2h_sdram0_READDATA_168,
	f2h_sdram0_READDATA_169,
	f2h_sdram0_READDATA_170,
	f2h_sdram0_READDATA_171,
	f2h_sdram0_READDATA_172,
	f2h_sdram0_READDATA_173,
	f2h_sdram0_READDATA_174,
	f2h_sdram0_READDATA_175,
	f2h_sdram0_READDATA_176,
	f2h_sdram0_READDATA_177,
	f2h_sdram0_READDATA_178,
	f2h_sdram0_READDATA_179,
	f2h_sdram0_READDATA_180,
	f2h_sdram0_READDATA_181,
	f2h_sdram0_READDATA_182,
	f2h_sdram0_READDATA_183,
	f2h_sdram0_READDATA_184,
	f2h_sdram0_READDATA_185,
	f2h_sdram0_READDATA_186,
	f2h_sdram0_READDATA_187,
	f2h_sdram0_READDATA_188,
	f2h_sdram0_READDATA_189,
	f2h_sdram0_READDATA_190,
	f2h_sdram0_READDATA_191,
	f2h_sdram0_READDATA_192,
	f2h_sdram0_READDATA_193,
	f2h_sdram0_READDATA_194,
	f2h_sdram0_READDATA_195,
	f2h_sdram0_READDATA_196,
	f2h_sdram0_READDATA_197,
	f2h_sdram0_READDATA_198,
	f2h_sdram0_READDATA_199,
	f2h_sdram0_READDATA_200,
	f2h_sdram0_READDATA_201,
	f2h_sdram0_READDATA_202,
	f2h_sdram0_READDATA_203,
	f2h_sdram0_READDATA_204,
	f2h_sdram0_READDATA_205,
	f2h_sdram0_READDATA_206,
	f2h_sdram0_READDATA_207,
	f2h_sdram0_READDATA_208,
	f2h_sdram0_READDATA_209,
	f2h_sdram0_READDATA_210,
	f2h_sdram0_READDATA_211,
	f2h_sdram0_READDATA_212,
	f2h_sdram0_READDATA_213,
	f2h_sdram0_READDATA_214,
	f2h_sdram0_READDATA_215,
	f2h_sdram0_READDATA_216,
	f2h_sdram0_READDATA_217,
	f2h_sdram0_READDATA_218,
	f2h_sdram0_READDATA_219,
	f2h_sdram0_READDATA_220,
	f2h_sdram0_READDATA_221,
	f2h_sdram0_READDATA_222,
	f2h_sdram0_READDATA_223,
	f2h_sdram0_READDATA_224,
	f2h_sdram0_READDATA_225,
	f2h_sdram0_READDATA_226,
	f2h_sdram0_READDATA_227,
	f2h_sdram0_READDATA_228,
	f2h_sdram0_READDATA_229,
	f2h_sdram0_READDATA_230,
	f2h_sdram0_READDATA_231,
	f2h_sdram0_READDATA_232,
	f2h_sdram0_READDATA_233,
	f2h_sdram0_READDATA_234,
	f2h_sdram0_READDATA_235,
	f2h_sdram0_READDATA_236,
	f2h_sdram0_READDATA_237,
	f2h_sdram0_READDATA_238,
	f2h_sdram0_READDATA_239,
	f2h_sdram0_READDATA_240,
	f2h_sdram0_READDATA_241,
	f2h_sdram0_READDATA_242,
	f2h_sdram0_READDATA_243,
	f2h_sdram0_READDATA_244,
	f2h_sdram0_READDATA_245,
	f2h_sdram0_READDATA_246,
	f2h_sdram0_READDATA_247,
	f2h_sdram0_READDATA_248,
	f2h_sdram0_READDATA_249,
	f2h_sdram0_READDATA_250,
	f2h_sdram0_READDATA_251,
	f2h_sdram0_READDATA_252,
	f2h_sdram0_READDATA_253,
	f2h_sdram0_READDATA_254,
	f2h_sdram0_READDATA_255,
	cmd_sink_ready,
	nonposted_cmd_accepted,
	WideOr1,
	src_payload_0,
	WideOr11,
	nonposted_cmd_accepted1,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_0,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	src_data_8,
	src_data_9,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_11,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	sdio_inst,
	intermediate_2,
	intermediate_3,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_10,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	intermediate_111,
	uart0_inst,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_f2h_stm_hw_events_stm_hwevents_0,
	hps_f2h_stm_hw_events_stm_hwevents_1,
	hps_f2h_stm_hw_events_stm_hwevents_2,
	hps_f2h_stm_hw_events_stm_hwevents_3,
	hps_f2h_stm_hw_events_stm_hwevents_4,
	hps_f2h_stm_hw_events_stm_hwevents_5,
	hps_f2h_stm_hw_events_stm_hwevents_6,
	hps_f2h_stm_hw_events_stm_hwevents_7,
	hps_f2h_stm_hw_events_stm_hwevents_8,
	hps_f2h_stm_hw_events_stm_hwevents_9,
	hps_f2h_stm_hw_events_stm_hwevents_10,
	hps_f2h_stm_hw_events_stm_hwevents_11,
	hps_f2h_stm_hw_events_stm_hwevents_12,
	hps_f2h_stm_hw_events_stm_hwevents_13,
	hps_f2h_stm_hw_events_stm_hwevents_14,
	hps_f2h_stm_hw_events_stm_hwevents_15,
	hps_f2h_stm_hw_events_stm_hwevents_16,
	hps_f2h_stm_hw_events_stm_hwevents_17,
	hps_f2h_stm_hw_events_stm_hwevents_18,
	hps_f2h_stm_hw_events_stm_hwevents_19,
	hps_f2h_stm_hw_events_stm_hwevents_20,
	hps_f2h_stm_hw_events_stm_hwevents_21,
	hps_f2h_stm_hw_events_stm_hwevents_22,
	hps_f2h_stm_hw_events_stm_hwevents_23,
	hps_f2h_stm_hw_events_stm_hwevents_24,
	hps_f2h_stm_hw_events_stm_hwevents_25,
	hps_f2h_stm_hw_events_stm_hwevents_26,
	hps_f2h_stm_hw_events_stm_hwevents_27,
	clk_clk,
	hps_hps_io_hps_io_emac1_inst_RXD0,
	hps_hps_io_hps_io_emac1_inst_RXD1,
	hps_hps_io_hps_io_emac1_inst_RXD2,
	hps_hps_io_hps_io_emac1_inst_RXD3,
	hps_hps_io_hps_io_emac1_inst_RX_CLK,
	hps_hps_io_hps_io_emac1_inst_RX_CTL,
	hps_hps_io_hps_io_uart0_inst_RX,
	memory_oct_rzqin,
	hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n,
	hps_f2h_sdram0_data_read,
	hps_f2h_sdram0_data_write,
	hps_f2h_sdram0_data_address_0,
	hps_f2h_sdram0_data_address_1,
	hps_f2h_sdram0_data_address_2,
	hps_f2h_sdram0_data_address_3,
	hps_f2h_sdram0_data_address_4,
	hps_f2h_sdram0_data_address_5,
	hps_f2h_sdram0_data_address_6,
	hps_f2h_sdram0_data_address_7,
	hps_f2h_sdram0_data_address_8,
	hps_f2h_sdram0_data_address_9,
	hps_f2h_sdram0_data_address_10,
	hps_f2h_sdram0_data_address_11,
	hps_f2h_sdram0_data_address_12,
	hps_f2h_sdram0_data_address_13,
	hps_f2h_sdram0_data_address_14,
	hps_f2h_sdram0_data_address_15,
	hps_f2h_sdram0_data_address_16,
	hps_f2h_sdram0_data_address_17,
	hps_f2h_sdram0_data_address_18,
	hps_f2h_sdram0_data_address_19,
	hps_f2h_sdram0_data_address_20,
	hps_f2h_sdram0_data_address_21,
	hps_f2h_sdram0_data_address_22,
	hps_f2h_sdram0_data_address_23,
	hps_f2h_sdram0_data_address_24,
	hps_f2h_sdram0_data_address_25,
	hps_f2h_sdram0_data_address_26,
	hps_f2h_sdram0_data_burstcount_0,
	hps_f2h_sdram0_data_burstcount_1,
	hps_f2h_sdram0_data_burstcount_2,
	hps_f2h_sdram0_data_burstcount_3,
	hps_f2h_sdram0_data_burstcount_4,
	hps_f2h_sdram0_data_burstcount_5,
	hps_f2h_sdram0_data_burstcount_6,
	hps_f2h_sdram0_data_burstcount_7,
	hps_f2h_sdram0_data_writedata_0,
	hps_f2h_sdram0_data_writedata_1,
	hps_f2h_sdram0_data_writedata_2,
	hps_f2h_sdram0_data_writedata_3,
	hps_f2h_sdram0_data_writedata_4,
	hps_f2h_sdram0_data_writedata_5,
	hps_f2h_sdram0_data_writedata_6,
	hps_f2h_sdram0_data_writedata_7,
	hps_f2h_sdram0_data_writedata_8,
	hps_f2h_sdram0_data_writedata_9,
	hps_f2h_sdram0_data_writedata_10,
	hps_f2h_sdram0_data_writedata_11,
	hps_f2h_sdram0_data_writedata_12,
	hps_f2h_sdram0_data_writedata_13,
	hps_f2h_sdram0_data_writedata_14,
	hps_f2h_sdram0_data_writedata_15,
	hps_f2h_sdram0_data_writedata_16,
	hps_f2h_sdram0_data_writedata_17,
	hps_f2h_sdram0_data_writedata_18,
	hps_f2h_sdram0_data_writedata_19,
	hps_f2h_sdram0_data_writedata_20,
	hps_f2h_sdram0_data_writedata_21,
	hps_f2h_sdram0_data_writedata_22,
	hps_f2h_sdram0_data_writedata_23,
	hps_f2h_sdram0_data_writedata_24,
	hps_f2h_sdram0_data_writedata_25,
	hps_f2h_sdram0_data_writedata_26,
	hps_f2h_sdram0_data_writedata_27,
	hps_f2h_sdram0_data_writedata_28,
	hps_f2h_sdram0_data_writedata_29,
	hps_f2h_sdram0_data_writedata_30,
	hps_f2h_sdram0_data_writedata_31,
	hps_f2h_sdram0_data_writedata_32,
	hps_f2h_sdram0_data_writedata_33,
	hps_f2h_sdram0_data_writedata_34,
	hps_f2h_sdram0_data_writedata_35,
	hps_f2h_sdram0_data_writedata_36,
	hps_f2h_sdram0_data_writedata_37,
	hps_f2h_sdram0_data_writedata_38,
	hps_f2h_sdram0_data_writedata_39,
	hps_f2h_sdram0_data_writedata_40,
	hps_f2h_sdram0_data_writedata_41,
	hps_f2h_sdram0_data_writedata_42,
	hps_f2h_sdram0_data_writedata_43,
	hps_f2h_sdram0_data_writedata_44,
	hps_f2h_sdram0_data_writedata_45,
	hps_f2h_sdram0_data_writedata_46,
	hps_f2h_sdram0_data_writedata_47,
	hps_f2h_sdram0_data_writedata_48,
	hps_f2h_sdram0_data_writedata_49,
	hps_f2h_sdram0_data_writedata_50,
	hps_f2h_sdram0_data_writedata_51,
	hps_f2h_sdram0_data_writedata_52,
	hps_f2h_sdram0_data_writedata_53,
	hps_f2h_sdram0_data_writedata_54,
	hps_f2h_sdram0_data_writedata_55,
	hps_f2h_sdram0_data_writedata_56,
	hps_f2h_sdram0_data_writedata_57,
	hps_f2h_sdram0_data_writedata_58,
	hps_f2h_sdram0_data_writedata_59,
	hps_f2h_sdram0_data_writedata_60,
	hps_f2h_sdram0_data_writedata_61,
	hps_f2h_sdram0_data_writedata_62,
	hps_f2h_sdram0_data_writedata_63,
	hps_f2h_sdram0_data_byteenable_0,
	hps_f2h_sdram0_data_byteenable_1,
	hps_f2h_sdram0_data_byteenable_2,
	hps_f2h_sdram0_data_byteenable_3,
	hps_f2h_sdram0_data_byteenable_4,
	hps_f2h_sdram0_data_byteenable_5,
	hps_f2h_sdram0_data_byteenable_6,
	hps_f2h_sdram0_data_byteenable_7,
	hps_f2h_sdram0_data_writedata_64,
	hps_f2h_sdram0_data_writedata_65,
	hps_f2h_sdram0_data_writedata_66,
	hps_f2h_sdram0_data_writedata_67,
	hps_f2h_sdram0_data_writedata_68,
	hps_f2h_sdram0_data_writedata_69,
	hps_f2h_sdram0_data_writedata_70,
	hps_f2h_sdram0_data_writedata_71,
	hps_f2h_sdram0_data_writedata_72,
	hps_f2h_sdram0_data_writedata_73,
	hps_f2h_sdram0_data_writedata_74,
	hps_f2h_sdram0_data_writedata_75,
	hps_f2h_sdram0_data_writedata_76,
	hps_f2h_sdram0_data_writedata_77,
	hps_f2h_sdram0_data_writedata_78,
	hps_f2h_sdram0_data_writedata_79,
	hps_f2h_sdram0_data_writedata_80,
	hps_f2h_sdram0_data_writedata_81,
	hps_f2h_sdram0_data_writedata_82,
	hps_f2h_sdram0_data_writedata_83,
	hps_f2h_sdram0_data_writedata_84,
	hps_f2h_sdram0_data_writedata_85,
	hps_f2h_sdram0_data_writedata_86,
	hps_f2h_sdram0_data_writedata_87,
	hps_f2h_sdram0_data_writedata_88,
	hps_f2h_sdram0_data_writedata_89,
	hps_f2h_sdram0_data_writedata_90,
	hps_f2h_sdram0_data_writedata_91,
	hps_f2h_sdram0_data_writedata_92,
	hps_f2h_sdram0_data_writedata_93,
	hps_f2h_sdram0_data_writedata_94,
	hps_f2h_sdram0_data_writedata_95,
	hps_f2h_sdram0_data_writedata_96,
	hps_f2h_sdram0_data_writedata_97,
	hps_f2h_sdram0_data_writedata_98,
	hps_f2h_sdram0_data_writedata_99,
	hps_f2h_sdram0_data_writedata_100,
	hps_f2h_sdram0_data_writedata_101,
	hps_f2h_sdram0_data_writedata_102,
	hps_f2h_sdram0_data_writedata_103,
	hps_f2h_sdram0_data_writedata_104,
	hps_f2h_sdram0_data_writedata_105,
	hps_f2h_sdram0_data_writedata_106,
	hps_f2h_sdram0_data_writedata_107,
	hps_f2h_sdram0_data_writedata_108,
	hps_f2h_sdram0_data_writedata_109,
	hps_f2h_sdram0_data_writedata_110,
	hps_f2h_sdram0_data_writedata_111,
	hps_f2h_sdram0_data_writedata_112,
	hps_f2h_sdram0_data_writedata_113,
	hps_f2h_sdram0_data_writedata_114,
	hps_f2h_sdram0_data_writedata_115,
	hps_f2h_sdram0_data_writedata_116,
	hps_f2h_sdram0_data_writedata_117,
	hps_f2h_sdram0_data_writedata_118,
	hps_f2h_sdram0_data_writedata_119,
	hps_f2h_sdram0_data_writedata_120,
	hps_f2h_sdram0_data_writedata_121,
	hps_f2h_sdram0_data_writedata_122,
	hps_f2h_sdram0_data_writedata_123,
	hps_f2h_sdram0_data_writedata_124,
	hps_f2h_sdram0_data_writedata_125,
	hps_f2h_sdram0_data_writedata_126,
	hps_f2h_sdram0_data_writedata_127,
	hps_f2h_sdram0_data_byteenable_8,
	hps_f2h_sdram0_data_byteenable_9,
	hps_f2h_sdram0_data_byteenable_10,
	hps_f2h_sdram0_data_byteenable_11,
	hps_f2h_sdram0_data_byteenable_12,
	hps_f2h_sdram0_data_byteenable_13,
	hps_f2h_sdram0_data_byteenable_14,
	hps_f2h_sdram0_data_byteenable_15,
	hps_f2h_sdram0_data_writedata_128,
	hps_f2h_sdram0_data_writedata_129,
	hps_f2h_sdram0_data_writedata_130,
	hps_f2h_sdram0_data_writedata_131,
	hps_f2h_sdram0_data_writedata_132,
	hps_f2h_sdram0_data_writedata_133,
	hps_f2h_sdram0_data_writedata_134,
	hps_f2h_sdram0_data_writedata_135,
	hps_f2h_sdram0_data_writedata_136,
	hps_f2h_sdram0_data_writedata_137,
	hps_f2h_sdram0_data_writedata_138,
	hps_f2h_sdram0_data_writedata_139,
	hps_f2h_sdram0_data_writedata_140,
	hps_f2h_sdram0_data_writedata_141,
	hps_f2h_sdram0_data_writedata_142,
	hps_f2h_sdram0_data_writedata_143,
	hps_f2h_sdram0_data_writedata_144,
	hps_f2h_sdram0_data_writedata_145,
	hps_f2h_sdram0_data_writedata_146,
	hps_f2h_sdram0_data_writedata_147,
	hps_f2h_sdram0_data_writedata_148,
	hps_f2h_sdram0_data_writedata_149,
	hps_f2h_sdram0_data_writedata_150,
	hps_f2h_sdram0_data_writedata_151,
	hps_f2h_sdram0_data_writedata_152,
	hps_f2h_sdram0_data_writedata_153,
	hps_f2h_sdram0_data_writedata_154,
	hps_f2h_sdram0_data_writedata_155,
	hps_f2h_sdram0_data_writedata_156,
	hps_f2h_sdram0_data_writedata_157,
	hps_f2h_sdram0_data_writedata_158,
	hps_f2h_sdram0_data_writedata_159,
	hps_f2h_sdram0_data_writedata_160,
	hps_f2h_sdram0_data_writedata_161,
	hps_f2h_sdram0_data_writedata_162,
	hps_f2h_sdram0_data_writedata_163,
	hps_f2h_sdram0_data_writedata_164,
	hps_f2h_sdram0_data_writedata_165,
	hps_f2h_sdram0_data_writedata_166,
	hps_f2h_sdram0_data_writedata_167,
	hps_f2h_sdram0_data_writedata_168,
	hps_f2h_sdram0_data_writedata_169,
	hps_f2h_sdram0_data_writedata_170,
	hps_f2h_sdram0_data_writedata_171,
	hps_f2h_sdram0_data_writedata_172,
	hps_f2h_sdram0_data_writedata_173,
	hps_f2h_sdram0_data_writedata_174,
	hps_f2h_sdram0_data_writedata_175,
	hps_f2h_sdram0_data_writedata_176,
	hps_f2h_sdram0_data_writedata_177,
	hps_f2h_sdram0_data_writedata_178,
	hps_f2h_sdram0_data_writedata_179,
	hps_f2h_sdram0_data_writedata_180,
	hps_f2h_sdram0_data_writedata_181,
	hps_f2h_sdram0_data_writedata_182,
	hps_f2h_sdram0_data_writedata_183,
	hps_f2h_sdram0_data_writedata_184,
	hps_f2h_sdram0_data_writedata_185,
	hps_f2h_sdram0_data_writedata_186,
	hps_f2h_sdram0_data_writedata_187,
	hps_f2h_sdram0_data_writedata_188,
	hps_f2h_sdram0_data_writedata_189,
	hps_f2h_sdram0_data_writedata_190,
	hps_f2h_sdram0_data_writedata_191,
	hps_f2h_sdram0_data_byteenable_16,
	hps_f2h_sdram0_data_byteenable_17,
	hps_f2h_sdram0_data_byteenable_18,
	hps_f2h_sdram0_data_byteenable_19,
	hps_f2h_sdram0_data_byteenable_20,
	hps_f2h_sdram0_data_byteenable_21,
	hps_f2h_sdram0_data_byteenable_22,
	hps_f2h_sdram0_data_byteenable_23,
	hps_f2h_sdram0_data_writedata_192,
	hps_f2h_sdram0_data_writedata_193,
	hps_f2h_sdram0_data_writedata_194,
	hps_f2h_sdram0_data_writedata_195,
	hps_f2h_sdram0_data_writedata_196,
	hps_f2h_sdram0_data_writedata_197,
	hps_f2h_sdram0_data_writedata_198,
	hps_f2h_sdram0_data_writedata_199,
	hps_f2h_sdram0_data_writedata_200,
	hps_f2h_sdram0_data_writedata_201,
	hps_f2h_sdram0_data_writedata_202,
	hps_f2h_sdram0_data_writedata_203,
	hps_f2h_sdram0_data_writedata_204,
	hps_f2h_sdram0_data_writedata_205,
	hps_f2h_sdram0_data_writedata_206,
	hps_f2h_sdram0_data_writedata_207,
	hps_f2h_sdram0_data_writedata_208,
	hps_f2h_sdram0_data_writedata_209,
	hps_f2h_sdram0_data_writedata_210,
	hps_f2h_sdram0_data_writedata_211,
	hps_f2h_sdram0_data_writedata_212,
	hps_f2h_sdram0_data_writedata_213,
	hps_f2h_sdram0_data_writedata_214,
	hps_f2h_sdram0_data_writedata_215,
	hps_f2h_sdram0_data_writedata_216,
	hps_f2h_sdram0_data_writedata_217,
	hps_f2h_sdram0_data_writedata_218,
	hps_f2h_sdram0_data_writedata_219,
	hps_f2h_sdram0_data_writedata_220,
	hps_f2h_sdram0_data_writedata_221,
	hps_f2h_sdram0_data_writedata_222,
	hps_f2h_sdram0_data_writedata_223,
	hps_f2h_sdram0_data_writedata_224,
	hps_f2h_sdram0_data_writedata_225,
	hps_f2h_sdram0_data_writedata_226,
	hps_f2h_sdram0_data_writedata_227,
	hps_f2h_sdram0_data_writedata_228,
	hps_f2h_sdram0_data_writedata_229,
	hps_f2h_sdram0_data_writedata_230,
	hps_f2h_sdram0_data_writedata_231,
	hps_f2h_sdram0_data_writedata_232,
	hps_f2h_sdram0_data_writedata_233,
	hps_f2h_sdram0_data_writedata_234,
	hps_f2h_sdram0_data_writedata_235,
	hps_f2h_sdram0_data_writedata_236,
	hps_f2h_sdram0_data_writedata_237,
	hps_f2h_sdram0_data_writedata_238,
	hps_f2h_sdram0_data_writedata_239,
	hps_f2h_sdram0_data_writedata_240,
	hps_f2h_sdram0_data_writedata_241,
	hps_f2h_sdram0_data_writedata_242,
	hps_f2h_sdram0_data_writedata_243,
	hps_f2h_sdram0_data_writedata_244,
	hps_f2h_sdram0_data_writedata_245,
	hps_f2h_sdram0_data_writedata_246,
	hps_f2h_sdram0_data_writedata_247,
	hps_f2h_sdram0_data_writedata_248,
	hps_f2h_sdram0_data_writedata_249,
	hps_f2h_sdram0_data_writedata_250,
	hps_f2h_sdram0_data_writedata_251,
	hps_f2h_sdram0_data_writedata_252,
	hps_f2h_sdram0_data_writedata_253,
	hps_f2h_sdram0_data_writedata_254,
	hps_f2h_sdram0_data_writedata_255,
	hps_f2h_sdram0_data_byteenable_24,
	hps_f2h_sdram0_data_byteenable_25,
	hps_f2h_sdram0_data_byteenable_26,
	hps_f2h_sdram0_data_byteenable_27,
	hps_f2h_sdram0_data_byteenable_28,
	hps_f2h_sdram0_data_byteenable_29,
	hps_f2h_sdram0_data_byteenable_30,
	hps_f2h_sdram0_data_byteenable_31)/* synthesis synthesis_greybox=0 */;
output 	h2f_cold_rst_n_0;
output 	h2f_pending_rst_req_n_0;
output 	h2f_rst_n_0;
output 	h2f_lw_ARVALID_0;
output 	h2f_lw_AWVALID_0;
output 	h2f_lw_BREADY_0;
output 	h2f_lw_RREADY_0;
output 	h2f_lw_WLAST_0;
output 	h2f_lw_WVALID_0;
output 	h2f_lw_ARADDR_0;
output 	h2f_lw_ARADDR_1;
output 	h2f_lw_ARADDR_2;
output 	h2f_lw_ARADDR_3;
output 	h2f_lw_ARADDR_4;
output 	h2f_lw_ARADDR_5;
output 	h2f_lw_ARADDR_6;
output 	h2f_lw_ARADDR_7;
output 	h2f_lw_ARADDR_8;
output 	h2f_lw_ARADDR_9;
output 	h2f_lw_ARADDR_10;
output 	h2f_lw_ARADDR_11;
output 	h2f_lw_ARADDR_12;
output 	h2f_lw_ARADDR_13;
output 	h2f_lw_ARADDR_14;
output 	h2f_lw_ARADDR_15;
output 	h2f_lw_ARADDR_16;
output 	h2f_lw_ARADDR_17;
output 	h2f_lw_ARADDR_18;
output 	h2f_lw_ARBURST_0;
output 	h2f_lw_ARBURST_1;
output 	h2f_lw_ARID_0;
output 	h2f_lw_ARID_1;
output 	h2f_lw_ARID_2;
output 	h2f_lw_ARID_3;
output 	h2f_lw_ARID_4;
output 	h2f_lw_ARID_5;
output 	h2f_lw_ARID_6;
output 	h2f_lw_ARID_7;
output 	h2f_lw_ARID_8;
output 	h2f_lw_ARID_9;
output 	h2f_lw_ARID_10;
output 	h2f_lw_ARID_11;
output 	h2f_lw_ARLEN_0;
output 	h2f_lw_ARLEN_1;
output 	h2f_lw_ARLEN_2;
output 	h2f_lw_ARLEN_3;
output 	h2f_lw_ARSIZE_0;
output 	h2f_lw_ARSIZE_1;
output 	h2f_lw_ARSIZE_2;
output 	h2f_lw_AWADDR_0;
output 	h2f_lw_AWADDR_1;
output 	h2f_lw_AWADDR_2;
output 	h2f_lw_AWADDR_3;
output 	h2f_lw_AWADDR_4;
output 	h2f_lw_AWADDR_5;
output 	h2f_lw_AWADDR_6;
output 	h2f_lw_AWADDR_7;
output 	h2f_lw_AWADDR_8;
output 	h2f_lw_AWADDR_9;
output 	h2f_lw_AWADDR_10;
output 	h2f_lw_AWADDR_11;
output 	h2f_lw_AWADDR_12;
output 	h2f_lw_AWADDR_13;
output 	h2f_lw_AWADDR_14;
output 	h2f_lw_AWADDR_15;
output 	h2f_lw_AWADDR_16;
output 	h2f_lw_AWADDR_17;
output 	h2f_lw_AWADDR_18;
output 	h2f_lw_AWBURST_0;
output 	h2f_lw_AWBURST_1;
output 	h2f_lw_AWID_0;
output 	h2f_lw_AWID_1;
output 	h2f_lw_AWID_2;
output 	h2f_lw_AWID_3;
output 	h2f_lw_AWID_4;
output 	h2f_lw_AWID_5;
output 	h2f_lw_AWID_6;
output 	h2f_lw_AWID_7;
output 	h2f_lw_AWID_8;
output 	h2f_lw_AWID_9;
output 	h2f_lw_AWID_10;
output 	h2f_lw_AWID_11;
output 	h2f_lw_AWLEN_0;
output 	h2f_lw_AWLEN_1;
output 	h2f_lw_AWLEN_2;
output 	h2f_lw_AWLEN_3;
output 	h2f_lw_AWSIZE_0;
output 	h2f_lw_AWSIZE_1;
output 	h2f_lw_AWSIZE_2;
output 	h2f_lw_WDATA_0;
output 	h2f_lw_WDATA_1;
output 	h2f_lw_WDATA_2;
output 	h2f_lw_WDATA_3;
output 	h2f_lw_WDATA_4;
output 	h2f_lw_WDATA_5;
output 	h2f_lw_WDATA_6;
output 	h2f_lw_WDATA_7;
output 	h2f_lw_WDATA_8;
output 	h2f_lw_WDATA_9;
output 	h2f_lw_WDATA_10;
output 	h2f_lw_WDATA_11;
output 	h2f_lw_WDATA_12;
output 	h2f_lw_WDATA_13;
output 	h2f_lw_WDATA_14;
output 	h2f_lw_WDATA_15;
output 	h2f_lw_WDATA_16;
output 	h2f_lw_WDATA_17;
output 	h2f_lw_WDATA_18;
output 	h2f_lw_WDATA_19;
output 	h2f_lw_WDATA_20;
output 	h2f_lw_WDATA_21;
output 	h2f_lw_WDATA_22;
output 	h2f_lw_WDATA_23;
output 	h2f_lw_WDATA_24;
output 	h2f_lw_WDATA_25;
output 	h2f_lw_WDATA_26;
output 	h2f_lw_WDATA_27;
output 	h2f_lw_WDATA_28;
output 	h2f_lw_WDATA_29;
output 	h2f_lw_WDATA_30;
output 	h2f_lw_WDATA_31;
output 	h2f_lw_WSTRB_0;
output 	h2f_lw_WSTRB_1;
output 	h2f_lw_WSTRB_2;
output 	h2f_lw_WSTRB_3;
output 	intermediate_1;
output 	f2h_sdram0_READDATAVALID_0;
output 	f2h_sdram0_READDATA_0;
output 	f2h_sdram0_READDATA_1;
output 	f2h_sdram0_READDATA_2;
output 	f2h_sdram0_READDATA_3;
output 	f2h_sdram0_READDATA_4;
output 	f2h_sdram0_READDATA_5;
output 	f2h_sdram0_READDATA_6;
output 	f2h_sdram0_READDATA_7;
output 	f2h_sdram0_READDATA_8;
output 	f2h_sdram0_READDATA_9;
output 	f2h_sdram0_READDATA_10;
output 	f2h_sdram0_READDATA_11;
output 	f2h_sdram0_READDATA_12;
output 	f2h_sdram0_READDATA_13;
output 	f2h_sdram0_READDATA_14;
output 	f2h_sdram0_READDATA_15;
output 	f2h_sdram0_READDATA_16;
output 	f2h_sdram0_READDATA_17;
output 	f2h_sdram0_READDATA_18;
output 	f2h_sdram0_READDATA_19;
output 	f2h_sdram0_READDATA_20;
output 	f2h_sdram0_READDATA_21;
output 	f2h_sdram0_READDATA_22;
output 	f2h_sdram0_READDATA_23;
output 	f2h_sdram0_READDATA_24;
output 	f2h_sdram0_READDATA_25;
output 	f2h_sdram0_READDATA_26;
output 	f2h_sdram0_READDATA_27;
output 	f2h_sdram0_READDATA_28;
output 	f2h_sdram0_READDATA_29;
output 	f2h_sdram0_READDATA_30;
output 	f2h_sdram0_READDATA_31;
output 	f2h_sdram0_READDATA_32;
output 	f2h_sdram0_READDATA_33;
output 	f2h_sdram0_READDATA_34;
output 	f2h_sdram0_READDATA_35;
output 	f2h_sdram0_READDATA_36;
output 	f2h_sdram0_READDATA_37;
output 	f2h_sdram0_READDATA_38;
output 	f2h_sdram0_READDATA_39;
output 	f2h_sdram0_READDATA_40;
output 	f2h_sdram0_READDATA_41;
output 	f2h_sdram0_READDATA_42;
output 	f2h_sdram0_READDATA_43;
output 	f2h_sdram0_READDATA_44;
output 	f2h_sdram0_READDATA_45;
output 	f2h_sdram0_READDATA_46;
output 	f2h_sdram0_READDATA_47;
output 	f2h_sdram0_READDATA_48;
output 	f2h_sdram0_READDATA_49;
output 	f2h_sdram0_READDATA_50;
output 	f2h_sdram0_READDATA_51;
output 	f2h_sdram0_READDATA_52;
output 	f2h_sdram0_READDATA_53;
output 	f2h_sdram0_READDATA_54;
output 	f2h_sdram0_READDATA_55;
output 	f2h_sdram0_READDATA_56;
output 	f2h_sdram0_READDATA_57;
output 	f2h_sdram0_READDATA_58;
output 	f2h_sdram0_READDATA_59;
output 	f2h_sdram0_READDATA_60;
output 	f2h_sdram0_READDATA_61;
output 	f2h_sdram0_READDATA_62;
output 	f2h_sdram0_READDATA_63;
output 	f2h_sdram0_READDATA_64;
output 	f2h_sdram0_READDATA_65;
output 	f2h_sdram0_READDATA_66;
output 	f2h_sdram0_READDATA_67;
output 	f2h_sdram0_READDATA_68;
output 	f2h_sdram0_READDATA_69;
output 	f2h_sdram0_READDATA_70;
output 	f2h_sdram0_READDATA_71;
output 	f2h_sdram0_READDATA_72;
output 	f2h_sdram0_READDATA_73;
output 	f2h_sdram0_READDATA_74;
output 	f2h_sdram0_READDATA_75;
output 	f2h_sdram0_READDATA_76;
output 	f2h_sdram0_READDATA_77;
output 	f2h_sdram0_READDATA_78;
output 	f2h_sdram0_READDATA_79;
output 	f2h_sdram0_READDATA_80;
output 	f2h_sdram0_READDATA_81;
output 	f2h_sdram0_READDATA_82;
output 	f2h_sdram0_READDATA_83;
output 	f2h_sdram0_READDATA_84;
output 	f2h_sdram0_READDATA_85;
output 	f2h_sdram0_READDATA_86;
output 	f2h_sdram0_READDATA_87;
output 	f2h_sdram0_READDATA_88;
output 	f2h_sdram0_READDATA_89;
output 	f2h_sdram0_READDATA_90;
output 	f2h_sdram0_READDATA_91;
output 	f2h_sdram0_READDATA_92;
output 	f2h_sdram0_READDATA_93;
output 	f2h_sdram0_READDATA_94;
output 	f2h_sdram0_READDATA_95;
output 	f2h_sdram0_READDATA_96;
output 	f2h_sdram0_READDATA_97;
output 	f2h_sdram0_READDATA_98;
output 	f2h_sdram0_READDATA_99;
output 	f2h_sdram0_READDATA_100;
output 	f2h_sdram0_READDATA_101;
output 	f2h_sdram0_READDATA_102;
output 	f2h_sdram0_READDATA_103;
output 	f2h_sdram0_READDATA_104;
output 	f2h_sdram0_READDATA_105;
output 	f2h_sdram0_READDATA_106;
output 	f2h_sdram0_READDATA_107;
output 	f2h_sdram0_READDATA_108;
output 	f2h_sdram0_READDATA_109;
output 	f2h_sdram0_READDATA_110;
output 	f2h_sdram0_READDATA_111;
output 	f2h_sdram0_READDATA_112;
output 	f2h_sdram0_READDATA_113;
output 	f2h_sdram0_READDATA_114;
output 	f2h_sdram0_READDATA_115;
output 	f2h_sdram0_READDATA_116;
output 	f2h_sdram0_READDATA_117;
output 	f2h_sdram0_READDATA_118;
output 	f2h_sdram0_READDATA_119;
output 	f2h_sdram0_READDATA_120;
output 	f2h_sdram0_READDATA_121;
output 	f2h_sdram0_READDATA_122;
output 	f2h_sdram0_READDATA_123;
output 	f2h_sdram0_READDATA_124;
output 	f2h_sdram0_READDATA_125;
output 	f2h_sdram0_READDATA_126;
output 	f2h_sdram0_READDATA_127;
output 	f2h_sdram0_READDATA_128;
output 	f2h_sdram0_READDATA_129;
output 	f2h_sdram0_READDATA_130;
output 	f2h_sdram0_READDATA_131;
output 	f2h_sdram0_READDATA_132;
output 	f2h_sdram0_READDATA_133;
output 	f2h_sdram0_READDATA_134;
output 	f2h_sdram0_READDATA_135;
output 	f2h_sdram0_READDATA_136;
output 	f2h_sdram0_READDATA_137;
output 	f2h_sdram0_READDATA_138;
output 	f2h_sdram0_READDATA_139;
output 	f2h_sdram0_READDATA_140;
output 	f2h_sdram0_READDATA_141;
output 	f2h_sdram0_READDATA_142;
output 	f2h_sdram0_READDATA_143;
output 	f2h_sdram0_READDATA_144;
output 	f2h_sdram0_READDATA_145;
output 	f2h_sdram0_READDATA_146;
output 	f2h_sdram0_READDATA_147;
output 	f2h_sdram0_READDATA_148;
output 	f2h_sdram0_READDATA_149;
output 	f2h_sdram0_READDATA_150;
output 	f2h_sdram0_READDATA_151;
output 	f2h_sdram0_READDATA_152;
output 	f2h_sdram0_READDATA_153;
output 	f2h_sdram0_READDATA_154;
output 	f2h_sdram0_READDATA_155;
output 	f2h_sdram0_READDATA_156;
output 	f2h_sdram0_READDATA_157;
output 	f2h_sdram0_READDATA_158;
output 	f2h_sdram0_READDATA_159;
output 	f2h_sdram0_READDATA_160;
output 	f2h_sdram0_READDATA_161;
output 	f2h_sdram0_READDATA_162;
output 	f2h_sdram0_READDATA_163;
output 	f2h_sdram0_READDATA_164;
output 	f2h_sdram0_READDATA_165;
output 	f2h_sdram0_READDATA_166;
output 	f2h_sdram0_READDATA_167;
output 	f2h_sdram0_READDATA_168;
output 	f2h_sdram0_READDATA_169;
output 	f2h_sdram0_READDATA_170;
output 	f2h_sdram0_READDATA_171;
output 	f2h_sdram0_READDATA_172;
output 	f2h_sdram0_READDATA_173;
output 	f2h_sdram0_READDATA_174;
output 	f2h_sdram0_READDATA_175;
output 	f2h_sdram0_READDATA_176;
output 	f2h_sdram0_READDATA_177;
output 	f2h_sdram0_READDATA_178;
output 	f2h_sdram0_READDATA_179;
output 	f2h_sdram0_READDATA_180;
output 	f2h_sdram0_READDATA_181;
output 	f2h_sdram0_READDATA_182;
output 	f2h_sdram0_READDATA_183;
output 	f2h_sdram0_READDATA_184;
output 	f2h_sdram0_READDATA_185;
output 	f2h_sdram0_READDATA_186;
output 	f2h_sdram0_READDATA_187;
output 	f2h_sdram0_READDATA_188;
output 	f2h_sdram0_READDATA_189;
output 	f2h_sdram0_READDATA_190;
output 	f2h_sdram0_READDATA_191;
output 	f2h_sdram0_READDATA_192;
output 	f2h_sdram0_READDATA_193;
output 	f2h_sdram0_READDATA_194;
output 	f2h_sdram0_READDATA_195;
output 	f2h_sdram0_READDATA_196;
output 	f2h_sdram0_READDATA_197;
output 	f2h_sdram0_READDATA_198;
output 	f2h_sdram0_READDATA_199;
output 	f2h_sdram0_READDATA_200;
output 	f2h_sdram0_READDATA_201;
output 	f2h_sdram0_READDATA_202;
output 	f2h_sdram0_READDATA_203;
output 	f2h_sdram0_READDATA_204;
output 	f2h_sdram0_READDATA_205;
output 	f2h_sdram0_READDATA_206;
output 	f2h_sdram0_READDATA_207;
output 	f2h_sdram0_READDATA_208;
output 	f2h_sdram0_READDATA_209;
output 	f2h_sdram0_READDATA_210;
output 	f2h_sdram0_READDATA_211;
output 	f2h_sdram0_READDATA_212;
output 	f2h_sdram0_READDATA_213;
output 	f2h_sdram0_READDATA_214;
output 	f2h_sdram0_READDATA_215;
output 	f2h_sdram0_READDATA_216;
output 	f2h_sdram0_READDATA_217;
output 	f2h_sdram0_READDATA_218;
output 	f2h_sdram0_READDATA_219;
output 	f2h_sdram0_READDATA_220;
output 	f2h_sdram0_READDATA_221;
output 	f2h_sdram0_READDATA_222;
output 	f2h_sdram0_READDATA_223;
output 	f2h_sdram0_READDATA_224;
output 	f2h_sdram0_READDATA_225;
output 	f2h_sdram0_READDATA_226;
output 	f2h_sdram0_READDATA_227;
output 	f2h_sdram0_READDATA_228;
output 	f2h_sdram0_READDATA_229;
output 	f2h_sdram0_READDATA_230;
output 	f2h_sdram0_READDATA_231;
output 	f2h_sdram0_READDATA_232;
output 	f2h_sdram0_READDATA_233;
output 	f2h_sdram0_READDATA_234;
output 	f2h_sdram0_READDATA_235;
output 	f2h_sdram0_READDATA_236;
output 	f2h_sdram0_READDATA_237;
output 	f2h_sdram0_READDATA_238;
output 	f2h_sdram0_READDATA_239;
output 	f2h_sdram0_READDATA_240;
output 	f2h_sdram0_READDATA_241;
output 	f2h_sdram0_READDATA_242;
output 	f2h_sdram0_READDATA_243;
output 	f2h_sdram0_READDATA_244;
output 	f2h_sdram0_READDATA_245;
output 	f2h_sdram0_READDATA_246;
output 	f2h_sdram0_READDATA_247;
output 	f2h_sdram0_READDATA_248;
output 	f2h_sdram0_READDATA_249;
output 	f2h_sdram0_READDATA_250;
output 	f2h_sdram0_READDATA_251;
output 	f2h_sdram0_READDATA_252;
output 	f2h_sdram0_READDATA_253;
output 	f2h_sdram0_READDATA_254;
output 	f2h_sdram0_READDATA_255;
input 	cmd_sink_ready;
input 	nonposted_cmd_accepted;
input 	WideOr1;
input 	src_payload_0;
input 	WideOr11;
input 	nonposted_cmd_accepted1;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_data_0;
input 	src_data_1;
input 	src_data_2;
input 	src_data_3;
input 	src_data_4;
input 	src_data_5;
input 	src_data_6;
input 	src_data_7;
input 	src_data_8;
input 	src_data_9;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	src_payload33;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_100;
input 	src_data_101;
input 	src_data_102;
input 	src_data_103;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_11;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	sdio_inst;
output 	intermediate_2;
output 	intermediate_3;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_10;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	intermediate_111;
output 	uart0_inst;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_f2h_stm_hw_events_stm_hwevents_0;
input 	hps_f2h_stm_hw_events_stm_hwevents_1;
input 	hps_f2h_stm_hw_events_stm_hwevents_2;
input 	hps_f2h_stm_hw_events_stm_hwevents_3;
input 	hps_f2h_stm_hw_events_stm_hwevents_4;
input 	hps_f2h_stm_hw_events_stm_hwevents_5;
input 	hps_f2h_stm_hw_events_stm_hwevents_6;
input 	hps_f2h_stm_hw_events_stm_hwevents_7;
input 	hps_f2h_stm_hw_events_stm_hwevents_8;
input 	hps_f2h_stm_hw_events_stm_hwevents_9;
input 	hps_f2h_stm_hw_events_stm_hwevents_10;
input 	hps_f2h_stm_hw_events_stm_hwevents_11;
input 	hps_f2h_stm_hw_events_stm_hwevents_12;
input 	hps_f2h_stm_hw_events_stm_hwevents_13;
input 	hps_f2h_stm_hw_events_stm_hwevents_14;
input 	hps_f2h_stm_hw_events_stm_hwevents_15;
input 	hps_f2h_stm_hw_events_stm_hwevents_16;
input 	hps_f2h_stm_hw_events_stm_hwevents_17;
input 	hps_f2h_stm_hw_events_stm_hwevents_18;
input 	hps_f2h_stm_hw_events_stm_hwevents_19;
input 	hps_f2h_stm_hw_events_stm_hwevents_20;
input 	hps_f2h_stm_hw_events_stm_hwevents_21;
input 	hps_f2h_stm_hw_events_stm_hwevents_22;
input 	hps_f2h_stm_hw_events_stm_hwevents_23;
input 	hps_f2h_stm_hw_events_stm_hwevents_24;
input 	hps_f2h_stm_hw_events_stm_hwevents_25;
input 	hps_f2h_stm_hw_events_stm_hwevents_26;
input 	hps_f2h_stm_hw_events_stm_hwevents_27;
input 	clk_clk;
input 	hps_hps_io_hps_io_emac1_inst_RXD0;
input 	hps_hps_io_hps_io_emac1_inst_RXD1;
input 	hps_hps_io_hps_io_emac1_inst_RXD2;
input 	hps_hps_io_hps_io_emac1_inst_RXD3;
input 	hps_hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_hps_io_hps_io_uart0_inst_RX;
input 	memory_oct_rzqin;
input 	hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n;
input 	hps_f2h_sdram0_data_read;
input 	hps_f2h_sdram0_data_write;
input 	hps_f2h_sdram0_data_address_0;
input 	hps_f2h_sdram0_data_address_1;
input 	hps_f2h_sdram0_data_address_2;
input 	hps_f2h_sdram0_data_address_3;
input 	hps_f2h_sdram0_data_address_4;
input 	hps_f2h_sdram0_data_address_5;
input 	hps_f2h_sdram0_data_address_6;
input 	hps_f2h_sdram0_data_address_7;
input 	hps_f2h_sdram0_data_address_8;
input 	hps_f2h_sdram0_data_address_9;
input 	hps_f2h_sdram0_data_address_10;
input 	hps_f2h_sdram0_data_address_11;
input 	hps_f2h_sdram0_data_address_12;
input 	hps_f2h_sdram0_data_address_13;
input 	hps_f2h_sdram0_data_address_14;
input 	hps_f2h_sdram0_data_address_15;
input 	hps_f2h_sdram0_data_address_16;
input 	hps_f2h_sdram0_data_address_17;
input 	hps_f2h_sdram0_data_address_18;
input 	hps_f2h_sdram0_data_address_19;
input 	hps_f2h_sdram0_data_address_20;
input 	hps_f2h_sdram0_data_address_21;
input 	hps_f2h_sdram0_data_address_22;
input 	hps_f2h_sdram0_data_address_23;
input 	hps_f2h_sdram0_data_address_24;
input 	hps_f2h_sdram0_data_address_25;
input 	hps_f2h_sdram0_data_address_26;
input 	hps_f2h_sdram0_data_burstcount_0;
input 	hps_f2h_sdram0_data_burstcount_1;
input 	hps_f2h_sdram0_data_burstcount_2;
input 	hps_f2h_sdram0_data_burstcount_3;
input 	hps_f2h_sdram0_data_burstcount_4;
input 	hps_f2h_sdram0_data_burstcount_5;
input 	hps_f2h_sdram0_data_burstcount_6;
input 	hps_f2h_sdram0_data_burstcount_7;
input 	hps_f2h_sdram0_data_writedata_0;
input 	hps_f2h_sdram0_data_writedata_1;
input 	hps_f2h_sdram0_data_writedata_2;
input 	hps_f2h_sdram0_data_writedata_3;
input 	hps_f2h_sdram0_data_writedata_4;
input 	hps_f2h_sdram0_data_writedata_5;
input 	hps_f2h_sdram0_data_writedata_6;
input 	hps_f2h_sdram0_data_writedata_7;
input 	hps_f2h_sdram0_data_writedata_8;
input 	hps_f2h_sdram0_data_writedata_9;
input 	hps_f2h_sdram0_data_writedata_10;
input 	hps_f2h_sdram0_data_writedata_11;
input 	hps_f2h_sdram0_data_writedata_12;
input 	hps_f2h_sdram0_data_writedata_13;
input 	hps_f2h_sdram0_data_writedata_14;
input 	hps_f2h_sdram0_data_writedata_15;
input 	hps_f2h_sdram0_data_writedata_16;
input 	hps_f2h_sdram0_data_writedata_17;
input 	hps_f2h_sdram0_data_writedata_18;
input 	hps_f2h_sdram0_data_writedata_19;
input 	hps_f2h_sdram0_data_writedata_20;
input 	hps_f2h_sdram0_data_writedata_21;
input 	hps_f2h_sdram0_data_writedata_22;
input 	hps_f2h_sdram0_data_writedata_23;
input 	hps_f2h_sdram0_data_writedata_24;
input 	hps_f2h_sdram0_data_writedata_25;
input 	hps_f2h_sdram0_data_writedata_26;
input 	hps_f2h_sdram0_data_writedata_27;
input 	hps_f2h_sdram0_data_writedata_28;
input 	hps_f2h_sdram0_data_writedata_29;
input 	hps_f2h_sdram0_data_writedata_30;
input 	hps_f2h_sdram0_data_writedata_31;
input 	hps_f2h_sdram0_data_writedata_32;
input 	hps_f2h_sdram0_data_writedata_33;
input 	hps_f2h_sdram0_data_writedata_34;
input 	hps_f2h_sdram0_data_writedata_35;
input 	hps_f2h_sdram0_data_writedata_36;
input 	hps_f2h_sdram0_data_writedata_37;
input 	hps_f2h_sdram0_data_writedata_38;
input 	hps_f2h_sdram0_data_writedata_39;
input 	hps_f2h_sdram0_data_writedata_40;
input 	hps_f2h_sdram0_data_writedata_41;
input 	hps_f2h_sdram0_data_writedata_42;
input 	hps_f2h_sdram0_data_writedata_43;
input 	hps_f2h_sdram0_data_writedata_44;
input 	hps_f2h_sdram0_data_writedata_45;
input 	hps_f2h_sdram0_data_writedata_46;
input 	hps_f2h_sdram0_data_writedata_47;
input 	hps_f2h_sdram0_data_writedata_48;
input 	hps_f2h_sdram0_data_writedata_49;
input 	hps_f2h_sdram0_data_writedata_50;
input 	hps_f2h_sdram0_data_writedata_51;
input 	hps_f2h_sdram0_data_writedata_52;
input 	hps_f2h_sdram0_data_writedata_53;
input 	hps_f2h_sdram0_data_writedata_54;
input 	hps_f2h_sdram0_data_writedata_55;
input 	hps_f2h_sdram0_data_writedata_56;
input 	hps_f2h_sdram0_data_writedata_57;
input 	hps_f2h_sdram0_data_writedata_58;
input 	hps_f2h_sdram0_data_writedata_59;
input 	hps_f2h_sdram0_data_writedata_60;
input 	hps_f2h_sdram0_data_writedata_61;
input 	hps_f2h_sdram0_data_writedata_62;
input 	hps_f2h_sdram0_data_writedata_63;
input 	hps_f2h_sdram0_data_byteenable_0;
input 	hps_f2h_sdram0_data_byteenable_1;
input 	hps_f2h_sdram0_data_byteenable_2;
input 	hps_f2h_sdram0_data_byteenable_3;
input 	hps_f2h_sdram0_data_byteenable_4;
input 	hps_f2h_sdram0_data_byteenable_5;
input 	hps_f2h_sdram0_data_byteenable_6;
input 	hps_f2h_sdram0_data_byteenable_7;
input 	hps_f2h_sdram0_data_writedata_64;
input 	hps_f2h_sdram0_data_writedata_65;
input 	hps_f2h_sdram0_data_writedata_66;
input 	hps_f2h_sdram0_data_writedata_67;
input 	hps_f2h_sdram0_data_writedata_68;
input 	hps_f2h_sdram0_data_writedata_69;
input 	hps_f2h_sdram0_data_writedata_70;
input 	hps_f2h_sdram0_data_writedata_71;
input 	hps_f2h_sdram0_data_writedata_72;
input 	hps_f2h_sdram0_data_writedata_73;
input 	hps_f2h_sdram0_data_writedata_74;
input 	hps_f2h_sdram0_data_writedata_75;
input 	hps_f2h_sdram0_data_writedata_76;
input 	hps_f2h_sdram0_data_writedata_77;
input 	hps_f2h_sdram0_data_writedata_78;
input 	hps_f2h_sdram0_data_writedata_79;
input 	hps_f2h_sdram0_data_writedata_80;
input 	hps_f2h_sdram0_data_writedata_81;
input 	hps_f2h_sdram0_data_writedata_82;
input 	hps_f2h_sdram0_data_writedata_83;
input 	hps_f2h_sdram0_data_writedata_84;
input 	hps_f2h_sdram0_data_writedata_85;
input 	hps_f2h_sdram0_data_writedata_86;
input 	hps_f2h_sdram0_data_writedata_87;
input 	hps_f2h_sdram0_data_writedata_88;
input 	hps_f2h_sdram0_data_writedata_89;
input 	hps_f2h_sdram0_data_writedata_90;
input 	hps_f2h_sdram0_data_writedata_91;
input 	hps_f2h_sdram0_data_writedata_92;
input 	hps_f2h_sdram0_data_writedata_93;
input 	hps_f2h_sdram0_data_writedata_94;
input 	hps_f2h_sdram0_data_writedata_95;
input 	hps_f2h_sdram0_data_writedata_96;
input 	hps_f2h_sdram0_data_writedata_97;
input 	hps_f2h_sdram0_data_writedata_98;
input 	hps_f2h_sdram0_data_writedata_99;
input 	hps_f2h_sdram0_data_writedata_100;
input 	hps_f2h_sdram0_data_writedata_101;
input 	hps_f2h_sdram0_data_writedata_102;
input 	hps_f2h_sdram0_data_writedata_103;
input 	hps_f2h_sdram0_data_writedata_104;
input 	hps_f2h_sdram0_data_writedata_105;
input 	hps_f2h_sdram0_data_writedata_106;
input 	hps_f2h_sdram0_data_writedata_107;
input 	hps_f2h_sdram0_data_writedata_108;
input 	hps_f2h_sdram0_data_writedata_109;
input 	hps_f2h_sdram0_data_writedata_110;
input 	hps_f2h_sdram0_data_writedata_111;
input 	hps_f2h_sdram0_data_writedata_112;
input 	hps_f2h_sdram0_data_writedata_113;
input 	hps_f2h_sdram0_data_writedata_114;
input 	hps_f2h_sdram0_data_writedata_115;
input 	hps_f2h_sdram0_data_writedata_116;
input 	hps_f2h_sdram0_data_writedata_117;
input 	hps_f2h_sdram0_data_writedata_118;
input 	hps_f2h_sdram0_data_writedata_119;
input 	hps_f2h_sdram0_data_writedata_120;
input 	hps_f2h_sdram0_data_writedata_121;
input 	hps_f2h_sdram0_data_writedata_122;
input 	hps_f2h_sdram0_data_writedata_123;
input 	hps_f2h_sdram0_data_writedata_124;
input 	hps_f2h_sdram0_data_writedata_125;
input 	hps_f2h_sdram0_data_writedata_126;
input 	hps_f2h_sdram0_data_writedata_127;
input 	hps_f2h_sdram0_data_byteenable_8;
input 	hps_f2h_sdram0_data_byteenable_9;
input 	hps_f2h_sdram0_data_byteenable_10;
input 	hps_f2h_sdram0_data_byteenable_11;
input 	hps_f2h_sdram0_data_byteenable_12;
input 	hps_f2h_sdram0_data_byteenable_13;
input 	hps_f2h_sdram0_data_byteenable_14;
input 	hps_f2h_sdram0_data_byteenable_15;
input 	hps_f2h_sdram0_data_writedata_128;
input 	hps_f2h_sdram0_data_writedata_129;
input 	hps_f2h_sdram0_data_writedata_130;
input 	hps_f2h_sdram0_data_writedata_131;
input 	hps_f2h_sdram0_data_writedata_132;
input 	hps_f2h_sdram0_data_writedata_133;
input 	hps_f2h_sdram0_data_writedata_134;
input 	hps_f2h_sdram0_data_writedata_135;
input 	hps_f2h_sdram0_data_writedata_136;
input 	hps_f2h_sdram0_data_writedata_137;
input 	hps_f2h_sdram0_data_writedata_138;
input 	hps_f2h_sdram0_data_writedata_139;
input 	hps_f2h_sdram0_data_writedata_140;
input 	hps_f2h_sdram0_data_writedata_141;
input 	hps_f2h_sdram0_data_writedata_142;
input 	hps_f2h_sdram0_data_writedata_143;
input 	hps_f2h_sdram0_data_writedata_144;
input 	hps_f2h_sdram0_data_writedata_145;
input 	hps_f2h_sdram0_data_writedata_146;
input 	hps_f2h_sdram0_data_writedata_147;
input 	hps_f2h_sdram0_data_writedata_148;
input 	hps_f2h_sdram0_data_writedata_149;
input 	hps_f2h_sdram0_data_writedata_150;
input 	hps_f2h_sdram0_data_writedata_151;
input 	hps_f2h_sdram0_data_writedata_152;
input 	hps_f2h_sdram0_data_writedata_153;
input 	hps_f2h_sdram0_data_writedata_154;
input 	hps_f2h_sdram0_data_writedata_155;
input 	hps_f2h_sdram0_data_writedata_156;
input 	hps_f2h_sdram0_data_writedata_157;
input 	hps_f2h_sdram0_data_writedata_158;
input 	hps_f2h_sdram0_data_writedata_159;
input 	hps_f2h_sdram0_data_writedata_160;
input 	hps_f2h_sdram0_data_writedata_161;
input 	hps_f2h_sdram0_data_writedata_162;
input 	hps_f2h_sdram0_data_writedata_163;
input 	hps_f2h_sdram0_data_writedata_164;
input 	hps_f2h_sdram0_data_writedata_165;
input 	hps_f2h_sdram0_data_writedata_166;
input 	hps_f2h_sdram0_data_writedata_167;
input 	hps_f2h_sdram0_data_writedata_168;
input 	hps_f2h_sdram0_data_writedata_169;
input 	hps_f2h_sdram0_data_writedata_170;
input 	hps_f2h_sdram0_data_writedata_171;
input 	hps_f2h_sdram0_data_writedata_172;
input 	hps_f2h_sdram0_data_writedata_173;
input 	hps_f2h_sdram0_data_writedata_174;
input 	hps_f2h_sdram0_data_writedata_175;
input 	hps_f2h_sdram0_data_writedata_176;
input 	hps_f2h_sdram0_data_writedata_177;
input 	hps_f2h_sdram0_data_writedata_178;
input 	hps_f2h_sdram0_data_writedata_179;
input 	hps_f2h_sdram0_data_writedata_180;
input 	hps_f2h_sdram0_data_writedata_181;
input 	hps_f2h_sdram0_data_writedata_182;
input 	hps_f2h_sdram0_data_writedata_183;
input 	hps_f2h_sdram0_data_writedata_184;
input 	hps_f2h_sdram0_data_writedata_185;
input 	hps_f2h_sdram0_data_writedata_186;
input 	hps_f2h_sdram0_data_writedata_187;
input 	hps_f2h_sdram0_data_writedata_188;
input 	hps_f2h_sdram0_data_writedata_189;
input 	hps_f2h_sdram0_data_writedata_190;
input 	hps_f2h_sdram0_data_writedata_191;
input 	hps_f2h_sdram0_data_byteenable_16;
input 	hps_f2h_sdram0_data_byteenable_17;
input 	hps_f2h_sdram0_data_byteenable_18;
input 	hps_f2h_sdram0_data_byteenable_19;
input 	hps_f2h_sdram0_data_byteenable_20;
input 	hps_f2h_sdram0_data_byteenable_21;
input 	hps_f2h_sdram0_data_byteenable_22;
input 	hps_f2h_sdram0_data_byteenable_23;
input 	hps_f2h_sdram0_data_writedata_192;
input 	hps_f2h_sdram0_data_writedata_193;
input 	hps_f2h_sdram0_data_writedata_194;
input 	hps_f2h_sdram0_data_writedata_195;
input 	hps_f2h_sdram0_data_writedata_196;
input 	hps_f2h_sdram0_data_writedata_197;
input 	hps_f2h_sdram0_data_writedata_198;
input 	hps_f2h_sdram0_data_writedata_199;
input 	hps_f2h_sdram0_data_writedata_200;
input 	hps_f2h_sdram0_data_writedata_201;
input 	hps_f2h_sdram0_data_writedata_202;
input 	hps_f2h_sdram0_data_writedata_203;
input 	hps_f2h_sdram0_data_writedata_204;
input 	hps_f2h_sdram0_data_writedata_205;
input 	hps_f2h_sdram0_data_writedata_206;
input 	hps_f2h_sdram0_data_writedata_207;
input 	hps_f2h_sdram0_data_writedata_208;
input 	hps_f2h_sdram0_data_writedata_209;
input 	hps_f2h_sdram0_data_writedata_210;
input 	hps_f2h_sdram0_data_writedata_211;
input 	hps_f2h_sdram0_data_writedata_212;
input 	hps_f2h_sdram0_data_writedata_213;
input 	hps_f2h_sdram0_data_writedata_214;
input 	hps_f2h_sdram0_data_writedata_215;
input 	hps_f2h_sdram0_data_writedata_216;
input 	hps_f2h_sdram0_data_writedata_217;
input 	hps_f2h_sdram0_data_writedata_218;
input 	hps_f2h_sdram0_data_writedata_219;
input 	hps_f2h_sdram0_data_writedata_220;
input 	hps_f2h_sdram0_data_writedata_221;
input 	hps_f2h_sdram0_data_writedata_222;
input 	hps_f2h_sdram0_data_writedata_223;
input 	hps_f2h_sdram0_data_writedata_224;
input 	hps_f2h_sdram0_data_writedata_225;
input 	hps_f2h_sdram0_data_writedata_226;
input 	hps_f2h_sdram0_data_writedata_227;
input 	hps_f2h_sdram0_data_writedata_228;
input 	hps_f2h_sdram0_data_writedata_229;
input 	hps_f2h_sdram0_data_writedata_230;
input 	hps_f2h_sdram0_data_writedata_231;
input 	hps_f2h_sdram0_data_writedata_232;
input 	hps_f2h_sdram0_data_writedata_233;
input 	hps_f2h_sdram0_data_writedata_234;
input 	hps_f2h_sdram0_data_writedata_235;
input 	hps_f2h_sdram0_data_writedata_236;
input 	hps_f2h_sdram0_data_writedata_237;
input 	hps_f2h_sdram0_data_writedata_238;
input 	hps_f2h_sdram0_data_writedata_239;
input 	hps_f2h_sdram0_data_writedata_240;
input 	hps_f2h_sdram0_data_writedata_241;
input 	hps_f2h_sdram0_data_writedata_242;
input 	hps_f2h_sdram0_data_writedata_243;
input 	hps_f2h_sdram0_data_writedata_244;
input 	hps_f2h_sdram0_data_writedata_245;
input 	hps_f2h_sdram0_data_writedata_246;
input 	hps_f2h_sdram0_data_writedata_247;
input 	hps_f2h_sdram0_data_writedata_248;
input 	hps_f2h_sdram0_data_writedata_249;
input 	hps_f2h_sdram0_data_writedata_250;
input 	hps_f2h_sdram0_data_writedata_251;
input 	hps_f2h_sdram0_data_writedata_252;
input 	hps_f2h_sdram0_data_writedata_253;
input 	hps_f2h_sdram0_data_writedata_254;
input 	hps_f2h_sdram0_data_writedata_255;
input 	hps_f2h_sdram0_data_byteenable_24;
input 	hps_f2h_sdram0_data_byteenable_25;
input 	hps_f2h_sdram0_data_byteenable_26;
input 	hps_f2h_sdram0_data_byteenable_27;
input 	hps_f2h_sdram0_data_byteenable_28;
input 	hps_f2h_sdram0_data_byteenable_29;
input 	hps_f2h_sdram0_data_byteenable_30;
input 	hps_f2h_sdram0_data_byteenable_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_terminal_qsys_hps_hps_io hps_io(
	.emac1_inst(emac1_inst),
	.emac1_inst1(emac1_inst1),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_11),
	.emac1_inst2(emac1_inst2),
	.emac1_inst3(emac1_inst3),
	.emac1_inst4(emac1_inst4),
	.emac1_inst5(emac1_inst5),
	.emac1_inst6(emac1_inst6),
	.sdio_inst(sdio_inst),
	.intermediate_2(intermediate_2),
	.intermediate_3(intermediate_3),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_10(intermediate_10),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.intermediate_11(intermediate_111),
	.uart0_inst(uart0_inst),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_hps_io_hps_io_emac1_inst_RXD0(hps_hps_io_hps_io_emac1_inst_RXD0),
	.hps_hps_io_hps_io_emac1_inst_RXD1(hps_hps_io_hps_io_emac1_inst_RXD1),
	.hps_hps_io_hps_io_emac1_inst_RXD2(hps_hps_io_hps_io_emac1_inst_RXD2),
	.hps_hps_io_hps_io_emac1_inst_RXD3(hps_hps_io_hps_io_emac1_inst_RXD3),
	.hps_hps_io_hps_io_emac1_inst_RX_CLK(hps_hps_io_hps_io_emac1_inst_RX_CLK),
	.hps_hps_io_hps_io_emac1_inst_RX_CTL(hps_hps_io_hps_io_emac1_inst_RX_CTL),
	.hps_hps_io_hps_io_uart0_inst_RX(hps_hps_io_hps_io_uart0_inst_RX),
	.memory_oct_rzqin(memory_oct_rzqin));

terminal_qsys_terminal_qsys_hps_fpga_interfaces fpga_interfaces(
	.h2f_cold_rst_n({h2f_cold_rst_n_0}),
	.h2f_pending_rst_req_n({h2f_pending_rst_req_n_0}),
	.h2f_rst_n({h2f_rst_n_0}),
	.h2f_lw_ARVALID({h2f_lw_ARVALID_0}),
	.h2f_lw_AWVALID({h2f_lw_AWVALID_0}),
	.h2f_lw_BREADY({h2f_lw_BREADY_0}),
	.h2f_lw_RREADY({h2f_lw_RREADY_0}),
	.h2f_lw_WLAST({h2f_lw_WLAST_0}),
	.h2f_lw_WVALID({h2f_lw_WVALID_0}),
	.h2f_lw_ARADDR({h2f_lw_ARADDR_unconnected_wire_20,h2f_lw_ARADDR_unconnected_wire_19,h2f_lw_ARADDR_18,h2f_lw_ARADDR_17,h2f_lw_ARADDR_16,h2f_lw_ARADDR_15,h2f_lw_ARADDR_14,h2f_lw_ARADDR_13,h2f_lw_ARADDR_12,h2f_lw_ARADDR_11,h2f_lw_ARADDR_10,h2f_lw_ARADDR_9,h2f_lw_ARADDR_8,h2f_lw_ARADDR_7,
h2f_lw_ARADDR_6,h2f_lw_ARADDR_5,h2f_lw_ARADDR_4,h2f_lw_ARADDR_3,h2f_lw_ARADDR_2,h2f_lw_ARADDR_1,h2f_lw_ARADDR_0}),
	.h2f_lw_ARBURST({h2f_lw_ARBURST_1,h2f_lw_ARBURST_0}),
	.h2f_lw_ARID({h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0}),
	.h2f_lw_ARLEN({h2f_lw_ARLEN_3,h2f_lw_ARLEN_2,h2f_lw_ARLEN_1,h2f_lw_ARLEN_0}),
	.h2f_lw_ARSIZE({h2f_lw_ARSIZE_2,h2f_lw_ARSIZE_1,h2f_lw_ARSIZE_0}),
	.h2f_lw_AWADDR({h2f_lw_AWADDR_unconnected_wire_20,h2f_lw_AWADDR_unconnected_wire_19,h2f_lw_AWADDR_18,h2f_lw_AWADDR_17,h2f_lw_AWADDR_16,h2f_lw_AWADDR_15,h2f_lw_AWADDR_14,h2f_lw_AWADDR_13,h2f_lw_AWADDR_12,h2f_lw_AWADDR_11,h2f_lw_AWADDR_10,h2f_lw_AWADDR_9,h2f_lw_AWADDR_8,h2f_lw_AWADDR_7,
h2f_lw_AWADDR_6,h2f_lw_AWADDR_5,h2f_lw_AWADDR_4,h2f_lw_AWADDR_3,h2f_lw_AWADDR_2,h2f_lw_AWADDR_1,h2f_lw_AWADDR_0}),
	.h2f_lw_AWBURST({h2f_lw_AWBURST_1,h2f_lw_AWBURST_0}),
	.h2f_lw_AWID({h2f_lw_AWID_11,h2f_lw_AWID_10,h2f_lw_AWID_9,h2f_lw_AWID_8,h2f_lw_AWID_7,h2f_lw_AWID_6,h2f_lw_AWID_5,h2f_lw_AWID_4,h2f_lw_AWID_3,h2f_lw_AWID_2,h2f_lw_AWID_1,h2f_lw_AWID_0}),
	.h2f_lw_AWLEN({h2f_lw_AWLEN_3,h2f_lw_AWLEN_2,h2f_lw_AWLEN_1,h2f_lw_AWLEN_0}),
	.h2f_lw_AWSIZE({h2f_lw_AWSIZE_2,h2f_lw_AWSIZE_1,h2f_lw_AWSIZE_0}),
	.h2f_lw_WDATA({h2f_lw_WDATA_31,h2f_lw_WDATA_30,h2f_lw_WDATA_29,h2f_lw_WDATA_28,h2f_lw_WDATA_27,h2f_lw_WDATA_26,h2f_lw_WDATA_25,h2f_lw_WDATA_24,h2f_lw_WDATA_23,h2f_lw_WDATA_22,h2f_lw_WDATA_21,h2f_lw_WDATA_20,h2f_lw_WDATA_19,h2f_lw_WDATA_18,h2f_lw_WDATA_17,h2f_lw_WDATA_16,h2f_lw_WDATA_15,
h2f_lw_WDATA_14,h2f_lw_WDATA_13,h2f_lw_WDATA_12,h2f_lw_WDATA_11,h2f_lw_WDATA_10,h2f_lw_WDATA_9,h2f_lw_WDATA_8,h2f_lw_WDATA_7,h2f_lw_WDATA_6,h2f_lw_WDATA_5,h2f_lw_WDATA_4,h2f_lw_WDATA_3,h2f_lw_WDATA_2,h2f_lw_WDATA_1,h2f_lw_WDATA_0}),
	.h2f_lw_WSTRB({h2f_lw_WSTRB_3,h2f_lw_WSTRB_2,h2f_lw_WSTRB_1,h2f_lw_WSTRB_0}),
	.f2h_sdram0_WAITREQUEST({intermediate_1}),
	.f2h_sdram0_READDATAVALID({f2h_sdram0_READDATAVALID_0}),
	.f2h_sdram0_READDATA({f2h_sdram0_READDATA_255,f2h_sdram0_READDATA_254,f2h_sdram0_READDATA_253,f2h_sdram0_READDATA_252,f2h_sdram0_READDATA_251,f2h_sdram0_READDATA_250,f2h_sdram0_READDATA_249,f2h_sdram0_READDATA_248,f2h_sdram0_READDATA_247,f2h_sdram0_READDATA_246,f2h_sdram0_READDATA_245,
f2h_sdram0_READDATA_244,f2h_sdram0_READDATA_243,f2h_sdram0_READDATA_242,f2h_sdram0_READDATA_241,f2h_sdram0_READDATA_240,f2h_sdram0_READDATA_239,f2h_sdram0_READDATA_238,f2h_sdram0_READDATA_237,f2h_sdram0_READDATA_236,f2h_sdram0_READDATA_235,f2h_sdram0_READDATA_234,
f2h_sdram0_READDATA_233,f2h_sdram0_READDATA_232,f2h_sdram0_READDATA_231,f2h_sdram0_READDATA_230,f2h_sdram0_READDATA_229,f2h_sdram0_READDATA_228,f2h_sdram0_READDATA_227,f2h_sdram0_READDATA_226,f2h_sdram0_READDATA_225,f2h_sdram0_READDATA_224,f2h_sdram0_READDATA_223,
f2h_sdram0_READDATA_222,f2h_sdram0_READDATA_221,f2h_sdram0_READDATA_220,f2h_sdram0_READDATA_219,f2h_sdram0_READDATA_218,f2h_sdram0_READDATA_217,f2h_sdram0_READDATA_216,f2h_sdram0_READDATA_215,f2h_sdram0_READDATA_214,f2h_sdram0_READDATA_213,f2h_sdram0_READDATA_212,
f2h_sdram0_READDATA_211,f2h_sdram0_READDATA_210,f2h_sdram0_READDATA_209,f2h_sdram0_READDATA_208,f2h_sdram0_READDATA_207,f2h_sdram0_READDATA_206,f2h_sdram0_READDATA_205,f2h_sdram0_READDATA_204,f2h_sdram0_READDATA_203,f2h_sdram0_READDATA_202,f2h_sdram0_READDATA_201,
f2h_sdram0_READDATA_200,f2h_sdram0_READDATA_199,f2h_sdram0_READDATA_198,f2h_sdram0_READDATA_197,f2h_sdram0_READDATA_196,f2h_sdram0_READDATA_195,f2h_sdram0_READDATA_194,f2h_sdram0_READDATA_193,f2h_sdram0_READDATA_192,f2h_sdram0_READDATA_191,f2h_sdram0_READDATA_190,
f2h_sdram0_READDATA_189,f2h_sdram0_READDATA_188,f2h_sdram0_READDATA_187,f2h_sdram0_READDATA_186,f2h_sdram0_READDATA_185,f2h_sdram0_READDATA_184,f2h_sdram0_READDATA_183,f2h_sdram0_READDATA_182,f2h_sdram0_READDATA_181,f2h_sdram0_READDATA_180,f2h_sdram0_READDATA_179,
f2h_sdram0_READDATA_178,f2h_sdram0_READDATA_177,f2h_sdram0_READDATA_176,f2h_sdram0_READDATA_175,f2h_sdram0_READDATA_174,f2h_sdram0_READDATA_173,f2h_sdram0_READDATA_172,f2h_sdram0_READDATA_171,f2h_sdram0_READDATA_170,f2h_sdram0_READDATA_169,f2h_sdram0_READDATA_168,
f2h_sdram0_READDATA_167,f2h_sdram0_READDATA_166,f2h_sdram0_READDATA_165,f2h_sdram0_READDATA_164,f2h_sdram0_READDATA_163,f2h_sdram0_READDATA_162,f2h_sdram0_READDATA_161,f2h_sdram0_READDATA_160,f2h_sdram0_READDATA_159,f2h_sdram0_READDATA_158,f2h_sdram0_READDATA_157,
f2h_sdram0_READDATA_156,f2h_sdram0_READDATA_155,f2h_sdram0_READDATA_154,f2h_sdram0_READDATA_153,f2h_sdram0_READDATA_152,f2h_sdram0_READDATA_151,f2h_sdram0_READDATA_150,f2h_sdram0_READDATA_149,f2h_sdram0_READDATA_148,f2h_sdram0_READDATA_147,f2h_sdram0_READDATA_146,
f2h_sdram0_READDATA_145,f2h_sdram0_READDATA_144,f2h_sdram0_READDATA_143,f2h_sdram0_READDATA_142,f2h_sdram0_READDATA_141,f2h_sdram0_READDATA_140,f2h_sdram0_READDATA_139,f2h_sdram0_READDATA_138,f2h_sdram0_READDATA_137,f2h_sdram0_READDATA_136,f2h_sdram0_READDATA_135,
f2h_sdram0_READDATA_134,f2h_sdram0_READDATA_133,f2h_sdram0_READDATA_132,f2h_sdram0_READDATA_131,f2h_sdram0_READDATA_130,f2h_sdram0_READDATA_129,f2h_sdram0_READDATA_128,f2h_sdram0_READDATA_127,f2h_sdram0_READDATA_126,f2h_sdram0_READDATA_125,f2h_sdram0_READDATA_124,
f2h_sdram0_READDATA_123,f2h_sdram0_READDATA_122,f2h_sdram0_READDATA_121,f2h_sdram0_READDATA_120,f2h_sdram0_READDATA_119,f2h_sdram0_READDATA_118,f2h_sdram0_READDATA_117,f2h_sdram0_READDATA_116,f2h_sdram0_READDATA_115,f2h_sdram0_READDATA_114,f2h_sdram0_READDATA_113,
f2h_sdram0_READDATA_112,f2h_sdram0_READDATA_111,f2h_sdram0_READDATA_110,f2h_sdram0_READDATA_109,f2h_sdram0_READDATA_108,f2h_sdram0_READDATA_107,f2h_sdram0_READDATA_106,f2h_sdram0_READDATA_105,f2h_sdram0_READDATA_104,f2h_sdram0_READDATA_103,f2h_sdram0_READDATA_102,
f2h_sdram0_READDATA_101,f2h_sdram0_READDATA_100,f2h_sdram0_READDATA_99,f2h_sdram0_READDATA_98,f2h_sdram0_READDATA_97,f2h_sdram0_READDATA_96,f2h_sdram0_READDATA_95,f2h_sdram0_READDATA_94,f2h_sdram0_READDATA_93,f2h_sdram0_READDATA_92,f2h_sdram0_READDATA_91,
f2h_sdram0_READDATA_90,f2h_sdram0_READDATA_89,f2h_sdram0_READDATA_88,f2h_sdram0_READDATA_87,f2h_sdram0_READDATA_86,f2h_sdram0_READDATA_85,f2h_sdram0_READDATA_84,f2h_sdram0_READDATA_83,f2h_sdram0_READDATA_82,f2h_sdram0_READDATA_81,f2h_sdram0_READDATA_80,
f2h_sdram0_READDATA_79,f2h_sdram0_READDATA_78,f2h_sdram0_READDATA_77,f2h_sdram0_READDATA_76,f2h_sdram0_READDATA_75,f2h_sdram0_READDATA_74,f2h_sdram0_READDATA_73,f2h_sdram0_READDATA_72,f2h_sdram0_READDATA_71,f2h_sdram0_READDATA_70,f2h_sdram0_READDATA_69,
f2h_sdram0_READDATA_68,f2h_sdram0_READDATA_67,f2h_sdram0_READDATA_66,f2h_sdram0_READDATA_65,f2h_sdram0_READDATA_64,f2h_sdram0_READDATA_63,f2h_sdram0_READDATA_62,f2h_sdram0_READDATA_61,f2h_sdram0_READDATA_60,f2h_sdram0_READDATA_59,f2h_sdram0_READDATA_58,
f2h_sdram0_READDATA_57,f2h_sdram0_READDATA_56,f2h_sdram0_READDATA_55,f2h_sdram0_READDATA_54,f2h_sdram0_READDATA_53,f2h_sdram0_READDATA_52,f2h_sdram0_READDATA_51,f2h_sdram0_READDATA_50,f2h_sdram0_READDATA_49,f2h_sdram0_READDATA_48,f2h_sdram0_READDATA_47,
f2h_sdram0_READDATA_46,f2h_sdram0_READDATA_45,f2h_sdram0_READDATA_44,f2h_sdram0_READDATA_43,f2h_sdram0_READDATA_42,f2h_sdram0_READDATA_41,f2h_sdram0_READDATA_40,f2h_sdram0_READDATA_39,f2h_sdram0_READDATA_38,f2h_sdram0_READDATA_37,f2h_sdram0_READDATA_36,
f2h_sdram0_READDATA_35,f2h_sdram0_READDATA_34,f2h_sdram0_READDATA_33,f2h_sdram0_READDATA_32,f2h_sdram0_READDATA_31,f2h_sdram0_READDATA_30,f2h_sdram0_READDATA_29,f2h_sdram0_READDATA_28,f2h_sdram0_READDATA_27,f2h_sdram0_READDATA_26,f2h_sdram0_READDATA_25,
f2h_sdram0_READDATA_24,f2h_sdram0_READDATA_23,f2h_sdram0_READDATA_22,f2h_sdram0_READDATA_21,f2h_sdram0_READDATA_20,f2h_sdram0_READDATA_19,f2h_sdram0_READDATA_18,f2h_sdram0_READDATA_17,f2h_sdram0_READDATA_16,f2h_sdram0_READDATA_15,f2h_sdram0_READDATA_14,
f2h_sdram0_READDATA_13,f2h_sdram0_READDATA_12,f2h_sdram0_READDATA_11,f2h_sdram0_READDATA_10,f2h_sdram0_READDATA_9,f2h_sdram0_READDATA_8,f2h_sdram0_READDATA_7,f2h_sdram0_READDATA_6,f2h_sdram0_READDATA_5,f2h_sdram0_READDATA_4,f2h_sdram0_READDATA_3,f2h_sdram0_READDATA_2,
f2h_sdram0_READDATA_1,f2h_sdram0_READDATA_0}),
	.h2f_lw_ARREADY({cmd_sink_ready}),
	.h2f_lw_AWREADY({nonposted_cmd_accepted}),
	.h2f_lw_BVALID({WideOr1}),
	.h2f_lw_RLAST({src_payload_0}),
	.h2f_lw_RVALID({WideOr11}),
	.h2f_lw_WREADY({nonposted_cmd_accepted1}),
	.h2f_lw_BID({src_payload11,src_payload10,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.h2f_lw_RDATA({src_payload33,src_payload32,src_payload31,src_payload30,src_payload29,src_payload28,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,
src_payload14,src_payload13,src_payload12,src_data_9,src_data_8,src_data_7,src_data_6,src_data_5,src_data_4,src_data_3,src_data_2,src_data_1,src_data_0}),
	.h2f_lw_RID({src_data_103,src_data_102,src_data_101,src_data_100,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92}),
	.f2h_stm_hwevents({hps_f2h_stm_hw_events_stm_hwevents_27,hps_f2h_stm_hw_events_stm_hwevents_26,hps_f2h_stm_hw_events_stm_hwevents_25,hps_f2h_stm_hw_events_stm_hwevents_24,hps_f2h_stm_hw_events_stm_hwevents_23,hps_f2h_stm_hw_events_stm_hwevents_22,
hps_f2h_stm_hw_events_stm_hwevents_21,hps_f2h_stm_hw_events_stm_hwevents_20,hps_f2h_stm_hw_events_stm_hwevents_19,hps_f2h_stm_hw_events_stm_hwevents_18,hps_f2h_stm_hw_events_stm_hwevents_17,hps_f2h_stm_hw_events_stm_hwevents_16,
hps_f2h_stm_hw_events_stm_hwevents_15,hps_f2h_stm_hw_events_stm_hwevents_14,hps_f2h_stm_hw_events_stm_hwevents_13,hps_f2h_stm_hw_events_stm_hwevents_12,hps_f2h_stm_hw_events_stm_hwevents_11,hps_f2h_stm_hw_events_stm_hwevents_10,
hps_f2h_stm_hw_events_stm_hwevents_9,hps_f2h_stm_hw_events_stm_hwevents_8,hps_f2h_stm_hw_events_stm_hwevents_7,hps_f2h_stm_hw_events_stm_hwevents_6,hps_f2h_stm_hw_events_stm_hwevents_5,hps_f2h_stm_hw_events_stm_hwevents_4,hps_f2h_stm_hw_events_stm_hwevents_3,
hps_f2h_stm_hw_events_stm_hwevents_2,hps_f2h_stm_hw_events_stm_hwevents_1,hps_f2h_stm_hw_events_stm_hwevents_0}),
	.h2f_lw_axi_clk({clk_clk}),
	.f2h_axi_clk({clk_clk}),
	.h2f_axi_clk({clk_clk}),
	.f2h_sdram0_clk({clk_clk}),
	.f2h_pending_rst_ack_n({hps_h2f_warm_reset_handshake_f2h_pending_rst_ack_n}),
	.f2h_sdram0_READ({hps_f2h_sdram0_data_read}),
	.f2h_sdram0_WRITE({hps_f2h_sdram0_data_write}),
	.f2h_sdram0_ADDRESS({hps_f2h_sdram0_data_address_26,hps_f2h_sdram0_data_address_25,hps_f2h_sdram0_data_address_24,hps_f2h_sdram0_data_address_23,hps_f2h_sdram0_data_address_22,hps_f2h_sdram0_data_address_21,hps_f2h_sdram0_data_address_20,hps_f2h_sdram0_data_address_19,
hps_f2h_sdram0_data_address_18,hps_f2h_sdram0_data_address_17,hps_f2h_sdram0_data_address_16,hps_f2h_sdram0_data_address_15,hps_f2h_sdram0_data_address_14,hps_f2h_sdram0_data_address_13,hps_f2h_sdram0_data_address_12,hps_f2h_sdram0_data_address_11,
hps_f2h_sdram0_data_address_10,hps_f2h_sdram0_data_address_9,hps_f2h_sdram0_data_address_8,hps_f2h_sdram0_data_address_7,hps_f2h_sdram0_data_address_6,hps_f2h_sdram0_data_address_5,hps_f2h_sdram0_data_address_4,hps_f2h_sdram0_data_address_3,
hps_f2h_sdram0_data_address_2,hps_f2h_sdram0_data_address_1,hps_f2h_sdram0_data_address_0}),
	.f2h_sdram0_BURSTCOUNT({hps_f2h_sdram0_data_burstcount_7,hps_f2h_sdram0_data_burstcount_6,hps_f2h_sdram0_data_burstcount_5,hps_f2h_sdram0_data_burstcount_4,hps_f2h_sdram0_data_burstcount_3,hps_f2h_sdram0_data_burstcount_2,hps_f2h_sdram0_data_burstcount_1,hps_f2h_sdram0_data_burstcount_0}),
	.f2h_sdram0_WRITEDATA({hps_f2h_sdram0_data_writedata_255,hps_f2h_sdram0_data_writedata_254,hps_f2h_sdram0_data_writedata_253,hps_f2h_sdram0_data_writedata_252,hps_f2h_sdram0_data_writedata_251,hps_f2h_sdram0_data_writedata_250,hps_f2h_sdram0_data_writedata_249,
hps_f2h_sdram0_data_writedata_248,hps_f2h_sdram0_data_writedata_247,hps_f2h_sdram0_data_writedata_246,hps_f2h_sdram0_data_writedata_245,hps_f2h_sdram0_data_writedata_244,hps_f2h_sdram0_data_writedata_243,hps_f2h_sdram0_data_writedata_242,
hps_f2h_sdram0_data_writedata_241,hps_f2h_sdram0_data_writedata_240,hps_f2h_sdram0_data_writedata_239,hps_f2h_sdram0_data_writedata_238,hps_f2h_sdram0_data_writedata_237,hps_f2h_sdram0_data_writedata_236,hps_f2h_sdram0_data_writedata_235,
hps_f2h_sdram0_data_writedata_234,hps_f2h_sdram0_data_writedata_233,hps_f2h_sdram0_data_writedata_232,hps_f2h_sdram0_data_writedata_231,hps_f2h_sdram0_data_writedata_230,hps_f2h_sdram0_data_writedata_229,hps_f2h_sdram0_data_writedata_228,
hps_f2h_sdram0_data_writedata_227,hps_f2h_sdram0_data_writedata_226,hps_f2h_sdram0_data_writedata_225,hps_f2h_sdram0_data_writedata_224,hps_f2h_sdram0_data_writedata_223,hps_f2h_sdram0_data_writedata_222,hps_f2h_sdram0_data_writedata_221,
hps_f2h_sdram0_data_writedata_220,hps_f2h_sdram0_data_writedata_219,hps_f2h_sdram0_data_writedata_218,hps_f2h_sdram0_data_writedata_217,hps_f2h_sdram0_data_writedata_216,hps_f2h_sdram0_data_writedata_215,hps_f2h_sdram0_data_writedata_214,
hps_f2h_sdram0_data_writedata_213,hps_f2h_sdram0_data_writedata_212,hps_f2h_sdram0_data_writedata_211,hps_f2h_sdram0_data_writedata_210,hps_f2h_sdram0_data_writedata_209,hps_f2h_sdram0_data_writedata_208,hps_f2h_sdram0_data_writedata_207,
hps_f2h_sdram0_data_writedata_206,hps_f2h_sdram0_data_writedata_205,hps_f2h_sdram0_data_writedata_204,hps_f2h_sdram0_data_writedata_203,hps_f2h_sdram0_data_writedata_202,hps_f2h_sdram0_data_writedata_201,hps_f2h_sdram0_data_writedata_200,
hps_f2h_sdram0_data_writedata_199,hps_f2h_sdram0_data_writedata_198,hps_f2h_sdram0_data_writedata_197,hps_f2h_sdram0_data_writedata_196,hps_f2h_sdram0_data_writedata_195,hps_f2h_sdram0_data_writedata_194,hps_f2h_sdram0_data_writedata_193,
hps_f2h_sdram0_data_writedata_192,hps_f2h_sdram0_data_writedata_191,hps_f2h_sdram0_data_writedata_190,hps_f2h_sdram0_data_writedata_189,hps_f2h_sdram0_data_writedata_188,hps_f2h_sdram0_data_writedata_187,hps_f2h_sdram0_data_writedata_186,
hps_f2h_sdram0_data_writedata_185,hps_f2h_sdram0_data_writedata_184,hps_f2h_sdram0_data_writedata_183,hps_f2h_sdram0_data_writedata_182,hps_f2h_sdram0_data_writedata_181,hps_f2h_sdram0_data_writedata_180,hps_f2h_sdram0_data_writedata_179,
hps_f2h_sdram0_data_writedata_178,hps_f2h_sdram0_data_writedata_177,hps_f2h_sdram0_data_writedata_176,hps_f2h_sdram0_data_writedata_175,hps_f2h_sdram0_data_writedata_174,hps_f2h_sdram0_data_writedata_173,hps_f2h_sdram0_data_writedata_172,
hps_f2h_sdram0_data_writedata_171,hps_f2h_sdram0_data_writedata_170,hps_f2h_sdram0_data_writedata_169,hps_f2h_sdram0_data_writedata_168,hps_f2h_sdram0_data_writedata_167,hps_f2h_sdram0_data_writedata_166,hps_f2h_sdram0_data_writedata_165,
hps_f2h_sdram0_data_writedata_164,hps_f2h_sdram0_data_writedata_163,hps_f2h_sdram0_data_writedata_162,hps_f2h_sdram0_data_writedata_161,hps_f2h_sdram0_data_writedata_160,hps_f2h_sdram0_data_writedata_159,hps_f2h_sdram0_data_writedata_158,
hps_f2h_sdram0_data_writedata_157,hps_f2h_sdram0_data_writedata_156,hps_f2h_sdram0_data_writedata_155,hps_f2h_sdram0_data_writedata_154,hps_f2h_sdram0_data_writedata_153,hps_f2h_sdram0_data_writedata_152,hps_f2h_sdram0_data_writedata_151,
hps_f2h_sdram0_data_writedata_150,hps_f2h_sdram0_data_writedata_149,hps_f2h_sdram0_data_writedata_148,hps_f2h_sdram0_data_writedata_147,hps_f2h_sdram0_data_writedata_146,hps_f2h_sdram0_data_writedata_145,hps_f2h_sdram0_data_writedata_144,
hps_f2h_sdram0_data_writedata_143,hps_f2h_sdram0_data_writedata_142,hps_f2h_sdram0_data_writedata_141,hps_f2h_sdram0_data_writedata_140,hps_f2h_sdram0_data_writedata_139,hps_f2h_sdram0_data_writedata_138,hps_f2h_sdram0_data_writedata_137,
hps_f2h_sdram0_data_writedata_136,hps_f2h_sdram0_data_writedata_135,hps_f2h_sdram0_data_writedata_134,hps_f2h_sdram0_data_writedata_133,hps_f2h_sdram0_data_writedata_132,hps_f2h_sdram0_data_writedata_131,hps_f2h_sdram0_data_writedata_130,
hps_f2h_sdram0_data_writedata_129,hps_f2h_sdram0_data_writedata_128,hps_f2h_sdram0_data_writedata_127,hps_f2h_sdram0_data_writedata_126,hps_f2h_sdram0_data_writedata_125,hps_f2h_sdram0_data_writedata_124,hps_f2h_sdram0_data_writedata_123,
hps_f2h_sdram0_data_writedata_122,hps_f2h_sdram0_data_writedata_121,hps_f2h_sdram0_data_writedata_120,hps_f2h_sdram0_data_writedata_119,hps_f2h_sdram0_data_writedata_118,hps_f2h_sdram0_data_writedata_117,hps_f2h_sdram0_data_writedata_116,
hps_f2h_sdram0_data_writedata_115,hps_f2h_sdram0_data_writedata_114,hps_f2h_sdram0_data_writedata_113,hps_f2h_sdram0_data_writedata_112,hps_f2h_sdram0_data_writedata_111,hps_f2h_sdram0_data_writedata_110,hps_f2h_sdram0_data_writedata_109,
hps_f2h_sdram0_data_writedata_108,hps_f2h_sdram0_data_writedata_107,hps_f2h_sdram0_data_writedata_106,hps_f2h_sdram0_data_writedata_105,hps_f2h_sdram0_data_writedata_104,hps_f2h_sdram0_data_writedata_103,hps_f2h_sdram0_data_writedata_102,
hps_f2h_sdram0_data_writedata_101,hps_f2h_sdram0_data_writedata_100,hps_f2h_sdram0_data_writedata_99,hps_f2h_sdram0_data_writedata_98,hps_f2h_sdram0_data_writedata_97,hps_f2h_sdram0_data_writedata_96,hps_f2h_sdram0_data_writedata_95,
hps_f2h_sdram0_data_writedata_94,hps_f2h_sdram0_data_writedata_93,hps_f2h_sdram0_data_writedata_92,hps_f2h_sdram0_data_writedata_91,hps_f2h_sdram0_data_writedata_90,hps_f2h_sdram0_data_writedata_89,hps_f2h_sdram0_data_writedata_88,hps_f2h_sdram0_data_writedata_87,
hps_f2h_sdram0_data_writedata_86,hps_f2h_sdram0_data_writedata_85,hps_f2h_sdram0_data_writedata_84,hps_f2h_sdram0_data_writedata_83,hps_f2h_sdram0_data_writedata_82,hps_f2h_sdram0_data_writedata_81,hps_f2h_sdram0_data_writedata_80,hps_f2h_sdram0_data_writedata_79,
hps_f2h_sdram0_data_writedata_78,hps_f2h_sdram0_data_writedata_77,hps_f2h_sdram0_data_writedata_76,hps_f2h_sdram0_data_writedata_75,hps_f2h_sdram0_data_writedata_74,hps_f2h_sdram0_data_writedata_73,hps_f2h_sdram0_data_writedata_72,hps_f2h_sdram0_data_writedata_71,
hps_f2h_sdram0_data_writedata_70,hps_f2h_sdram0_data_writedata_69,hps_f2h_sdram0_data_writedata_68,hps_f2h_sdram0_data_writedata_67,hps_f2h_sdram0_data_writedata_66,hps_f2h_sdram0_data_writedata_65,hps_f2h_sdram0_data_writedata_64,hps_f2h_sdram0_data_writedata_63,
hps_f2h_sdram0_data_writedata_62,hps_f2h_sdram0_data_writedata_61,hps_f2h_sdram0_data_writedata_60,hps_f2h_sdram0_data_writedata_59,hps_f2h_sdram0_data_writedata_58,hps_f2h_sdram0_data_writedata_57,hps_f2h_sdram0_data_writedata_56,hps_f2h_sdram0_data_writedata_55,
hps_f2h_sdram0_data_writedata_54,hps_f2h_sdram0_data_writedata_53,hps_f2h_sdram0_data_writedata_52,hps_f2h_sdram0_data_writedata_51,hps_f2h_sdram0_data_writedata_50,hps_f2h_sdram0_data_writedata_49,hps_f2h_sdram0_data_writedata_48,hps_f2h_sdram0_data_writedata_47,
hps_f2h_sdram0_data_writedata_46,hps_f2h_sdram0_data_writedata_45,hps_f2h_sdram0_data_writedata_44,hps_f2h_sdram0_data_writedata_43,hps_f2h_sdram0_data_writedata_42,hps_f2h_sdram0_data_writedata_41,hps_f2h_sdram0_data_writedata_40,hps_f2h_sdram0_data_writedata_39,
hps_f2h_sdram0_data_writedata_38,hps_f2h_sdram0_data_writedata_37,hps_f2h_sdram0_data_writedata_36,hps_f2h_sdram0_data_writedata_35,hps_f2h_sdram0_data_writedata_34,hps_f2h_sdram0_data_writedata_33,hps_f2h_sdram0_data_writedata_32,hps_f2h_sdram0_data_writedata_31,
hps_f2h_sdram0_data_writedata_30,hps_f2h_sdram0_data_writedata_29,hps_f2h_sdram0_data_writedata_28,hps_f2h_sdram0_data_writedata_27,hps_f2h_sdram0_data_writedata_26,hps_f2h_sdram0_data_writedata_25,hps_f2h_sdram0_data_writedata_24,hps_f2h_sdram0_data_writedata_23,
hps_f2h_sdram0_data_writedata_22,hps_f2h_sdram0_data_writedata_21,hps_f2h_sdram0_data_writedata_20,hps_f2h_sdram0_data_writedata_19,hps_f2h_sdram0_data_writedata_18,hps_f2h_sdram0_data_writedata_17,hps_f2h_sdram0_data_writedata_16,hps_f2h_sdram0_data_writedata_15,
hps_f2h_sdram0_data_writedata_14,hps_f2h_sdram0_data_writedata_13,hps_f2h_sdram0_data_writedata_12,hps_f2h_sdram0_data_writedata_11,hps_f2h_sdram0_data_writedata_10,hps_f2h_sdram0_data_writedata_9,hps_f2h_sdram0_data_writedata_8,hps_f2h_sdram0_data_writedata_7,
hps_f2h_sdram0_data_writedata_6,hps_f2h_sdram0_data_writedata_5,hps_f2h_sdram0_data_writedata_4,hps_f2h_sdram0_data_writedata_3,hps_f2h_sdram0_data_writedata_2,hps_f2h_sdram0_data_writedata_1,hps_f2h_sdram0_data_writedata_0}),
	.f2h_sdram0_BYTEENABLE({hps_f2h_sdram0_data_byteenable_31,hps_f2h_sdram0_data_byteenable_30,hps_f2h_sdram0_data_byteenable_29,hps_f2h_sdram0_data_byteenable_28,hps_f2h_sdram0_data_byteenable_27,hps_f2h_sdram0_data_byteenable_26,hps_f2h_sdram0_data_byteenable_25,
hps_f2h_sdram0_data_byteenable_24,hps_f2h_sdram0_data_byteenable_23,hps_f2h_sdram0_data_byteenable_22,hps_f2h_sdram0_data_byteenable_21,hps_f2h_sdram0_data_byteenable_20,hps_f2h_sdram0_data_byteenable_19,hps_f2h_sdram0_data_byteenable_18,
hps_f2h_sdram0_data_byteenable_17,hps_f2h_sdram0_data_byteenable_16,hps_f2h_sdram0_data_byteenable_15,hps_f2h_sdram0_data_byteenable_14,hps_f2h_sdram0_data_byteenable_13,hps_f2h_sdram0_data_byteenable_12,hps_f2h_sdram0_data_byteenable_11,
hps_f2h_sdram0_data_byteenable_10,hps_f2h_sdram0_data_byteenable_9,hps_f2h_sdram0_data_byteenable_8,hps_f2h_sdram0_data_byteenable_7,hps_f2h_sdram0_data_byteenable_6,hps_f2h_sdram0_data_byteenable_5,hps_f2h_sdram0_data_byteenable_4,
hps_f2h_sdram0_data_byteenable_3,hps_f2h_sdram0_data_byteenable_2,hps_f2h_sdram0_data_byteenable_1,hps_f2h_sdram0_data_byteenable_0}));

endmodule

module terminal_qsys_terminal_qsys_hps_fpga_interfaces (
	h2f_cold_rst_n,
	h2f_pending_rst_req_n,
	h2f_rst_n,
	h2f_lw_ARVALID,
	h2f_lw_AWVALID,
	h2f_lw_BREADY,
	h2f_lw_RREADY,
	h2f_lw_WLAST,
	h2f_lw_WVALID,
	h2f_lw_ARADDR,
	h2f_lw_ARBURST,
	h2f_lw_ARID,
	h2f_lw_ARLEN,
	h2f_lw_ARSIZE,
	h2f_lw_AWADDR,
	h2f_lw_AWBURST,
	h2f_lw_AWID,
	h2f_lw_AWLEN,
	h2f_lw_AWSIZE,
	h2f_lw_WDATA,
	h2f_lw_WSTRB,
	f2h_sdram0_WAITREQUEST,
	f2h_sdram0_READDATAVALID,
	f2h_sdram0_READDATA,
	h2f_lw_ARREADY,
	h2f_lw_AWREADY,
	h2f_lw_BVALID,
	h2f_lw_RLAST,
	h2f_lw_RVALID,
	h2f_lw_WREADY,
	h2f_lw_BID,
	h2f_lw_RDATA,
	h2f_lw_RID,
	f2h_stm_hwevents,
	h2f_lw_axi_clk,
	f2h_axi_clk,
	h2f_axi_clk,
	f2h_sdram0_clk,
	f2h_pending_rst_ack_n,
	f2h_sdram0_READ,
	f2h_sdram0_WRITE,
	f2h_sdram0_ADDRESS,
	f2h_sdram0_BURSTCOUNT,
	f2h_sdram0_WRITEDATA,
	f2h_sdram0_BYTEENABLE)/* synthesis synthesis_greybox=0 */;
output 	[0:0] h2f_cold_rst_n;
output 	[0:0] h2f_pending_rst_req_n;
output 	[0:0] h2f_rst_n;
output 	[0:0] h2f_lw_ARVALID;
output 	[0:0] h2f_lw_AWVALID;
output 	[0:0] h2f_lw_BREADY;
output 	[0:0] h2f_lw_RREADY;
output 	[0:0] h2f_lw_WLAST;
output 	[0:0] h2f_lw_WVALID;
output 	[20:0] h2f_lw_ARADDR;
output 	[1:0] h2f_lw_ARBURST;
output 	[11:0] h2f_lw_ARID;
output 	[3:0] h2f_lw_ARLEN;
output 	[2:0] h2f_lw_ARSIZE;
output 	[20:0] h2f_lw_AWADDR;
output 	[1:0] h2f_lw_AWBURST;
output 	[11:0] h2f_lw_AWID;
output 	[3:0] h2f_lw_AWLEN;
output 	[2:0] h2f_lw_AWSIZE;
output 	[31:0] h2f_lw_WDATA;
output 	[3:0] h2f_lw_WSTRB;
output 	[0:0] f2h_sdram0_WAITREQUEST;
output 	[0:0] f2h_sdram0_READDATAVALID;
output 	[255:0] f2h_sdram0_READDATA;
input 	[0:0] h2f_lw_ARREADY;
input 	[0:0] h2f_lw_AWREADY;
input 	[0:0] h2f_lw_BVALID;
input 	[0:0] h2f_lw_RLAST;
input 	[0:0] h2f_lw_RVALID;
input 	[0:0] h2f_lw_WREADY;
input 	[11:0] h2f_lw_BID;
input 	[31:0] h2f_lw_RDATA;
input 	[11:0] h2f_lw_RID;
input 	[27:0] f2h_stm_hwevents;
input 	[0:0] h2f_lw_axi_clk;
input 	[0:0] f2h_axi_clk;
input 	[0:0] h2f_axi_clk;
input 	[0:0] f2h_sdram0_clk;
input 	[0:0] f2h_pending_rst_ack_n;
input 	[0:0] f2h_sdram0_READ;
input 	[0:0] f2h_sdram0_WRITE;
input 	[26:0] f2h_sdram0_ADDRESS;
input 	[7:0] f2h_sdram0_BURSTCOUNT;
input 	[255:0] f2h_sdram0_WRITEDATA;
input 	[31:0] f2h_sdram0_BYTEENABLE;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \debug_apb~O_P_ADDR_31 ;
wire \stm_event~fake_dout ;
wire \tpiu~trace_data ;
wire \tpiu~O_TRACE_DATA1 ;
wire \tpiu~O_TRACE_DATA2 ;
wire \tpiu~O_TRACE_DATA3 ;
wire \tpiu~O_TRACE_DATA4 ;
wire \tpiu~O_TRACE_DATA5 ;
wire \tpiu~O_TRACE_DATA6 ;
wire \tpiu~O_TRACE_DATA7 ;
wire \tpiu~O_TRACE_DATA8 ;
wire \tpiu~O_TRACE_DATA9 ;
wire \tpiu~O_TRACE_DATA10 ;
wire \tpiu~O_TRACE_DATA11 ;
wire \tpiu~O_TRACE_DATA12 ;
wire \tpiu~O_TRACE_DATA13 ;
wire \tpiu~O_TRACE_DATA14 ;
wire \tpiu~O_TRACE_DATA15 ;
wire \tpiu~O_TRACE_DATA16 ;
wire \tpiu~O_TRACE_DATA17 ;
wire \tpiu~O_TRACE_DATA18 ;
wire \tpiu~O_TRACE_DATA19 ;
wire \tpiu~O_TRACE_DATA20 ;
wire \tpiu~O_TRACE_DATA21 ;
wire \tpiu~O_TRACE_DATA22 ;
wire \tpiu~O_TRACE_DATA23 ;
wire \tpiu~O_TRACE_DATA24 ;
wire \tpiu~O_TRACE_DATA25 ;
wire \tpiu~O_TRACE_DATA26 ;
wire \tpiu~O_TRACE_DATA27 ;
wire \tpiu~O_TRACE_DATA28 ;
wire \tpiu~O_TRACE_DATA29 ;
wire \tpiu~O_TRACE_DATA30 ;
wire \tpiu~O_TRACE_DATA31 ;
wire \boot_from_fpga~fake_dout ;
wire \f2h_ARREADY[0] ;
wire \h2f_ARADDR[0] ;
wire \h2f_ARADDR[1] ;
wire \h2f_ARADDR[2] ;
wire \h2f_ARADDR[3] ;
wire \h2f_ARADDR[4] ;
wire \h2f_ARADDR[5] ;
wire \h2f_ARADDR[6] ;
wire \h2f_ARADDR[7] ;
wire \h2f_ARADDR[8] ;
wire \h2f_ARADDR[9] ;
wire \h2f_ARADDR[10] ;
wire \h2f_ARADDR[11] ;
wire \h2f_ARADDR[12] ;
wire \h2f_ARADDR[13] ;
wire \h2f_ARADDR[14] ;
wire \h2f_ARADDR[15] ;
wire \h2f_ARADDR[16] ;
wire \h2f_ARADDR[17] ;
wire \h2f_ARADDR[18] ;
wire \h2f_ARADDR[19] ;
wire \h2f_ARADDR[20] ;
wire \h2f_ARADDR[21] ;
wire \h2f_ARADDR[22] ;
wire \h2f_ARADDR[23] ;
wire \h2f_ARADDR[24] ;
wire \h2f_ARADDR[25] ;
wire \h2f_ARADDR[26] ;
wire \h2f_ARADDR[27] ;
wire \h2f_ARADDR[28] ;
wire \h2f_ARADDR[29] ;
wire \h2f_lw_ARADDR[19] ;
wire \h2f_lw_ARADDR[20] ;
wire \f2sdram~O_BONDING_OUT_10 ;
wire \f2sdram~O_BONDING_OUT_11 ;
wire \f2sdram~O_BONDING_OUT_12 ;
wire \f2sdram~O_BONDING_OUT_13 ;
wire \intermediate[12]~combout ;

wire [31:0] tpiu_TRACE_DATA_bus;
wire [29:0] hps2fpga_ARADDR_bus;
wire [20:0] hps2fpga_light_weight_ARADDR_bus;
wire [1:0] hps2fpga_light_weight_ARBURST_bus;
wire [11:0] hps2fpga_light_weight_ARID_bus;
wire [3:0] hps2fpga_light_weight_ARLEN_bus;
wire [2:0] hps2fpga_light_weight_ARSIZE_bus;
wire [20:0] hps2fpga_light_weight_AWADDR_bus;
wire [1:0] hps2fpga_light_weight_AWBURST_bus;
wire [11:0] hps2fpga_light_weight_AWID_bus;
wire [3:0] hps2fpga_light_weight_AWLEN_bus;
wire [2:0] hps2fpga_light_weight_AWSIZE_bus;
wire [31:0] hps2fpga_light_weight_WDATA_bus;
wire [3:0] hps2fpga_light_weight_WSTRB_bus;
wire [3:0] f2sdram_BONDING_OUT_1_bus;
wire [79:0] f2sdram_RD_DATA_0_bus;
wire [79:0] f2sdram_RD_DATA_1_bus;
wire [79:0] f2sdram_RD_DATA_2_bus;
wire [79:0] f2sdram_RD_DATA_3_bus;

assign \tpiu~trace_data  = tpiu_TRACE_DATA_bus[0];
assign \tpiu~O_TRACE_DATA1  = tpiu_TRACE_DATA_bus[1];
assign \tpiu~O_TRACE_DATA2  = tpiu_TRACE_DATA_bus[2];
assign \tpiu~O_TRACE_DATA3  = tpiu_TRACE_DATA_bus[3];
assign \tpiu~O_TRACE_DATA4  = tpiu_TRACE_DATA_bus[4];
assign \tpiu~O_TRACE_DATA5  = tpiu_TRACE_DATA_bus[5];
assign \tpiu~O_TRACE_DATA6  = tpiu_TRACE_DATA_bus[6];
assign \tpiu~O_TRACE_DATA7  = tpiu_TRACE_DATA_bus[7];
assign \tpiu~O_TRACE_DATA8  = tpiu_TRACE_DATA_bus[8];
assign \tpiu~O_TRACE_DATA9  = tpiu_TRACE_DATA_bus[9];
assign \tpiu~O_TRACE_DATA10  = tpiu_TRACE_DATA_bus[10];
assign \tpiu~O_TRACE_DATA11  = tpiu_TRACE_DATA_bus[11];
assign \tpiu~O_TRACE_DATA12  = tpiu_TRACE_DATA_bus[12];
assign \tpiu~O_TRACE_DATA13  = tpiu_TRACE_DATA_bus[13];
assign \tpiu~O_TRACE_DATA14  = tpiu_TRACE_DATA_bus[14];
assign \tpiu~O_TRACE_DATA15  = tpiu_TRACE_DATA_bus[15];
assign \tpiu~O_TRACE_DATA16  = tpiu_TRACE_DATA_bus[16];
assign \tpiu~O_TRACE_DATA17  = tpiu_TRACE_DATA_bus[17];
assign \tpiu~O_TRACE_DATA18  = tpiu_TRACE_DATA_bus[18];
assign \tpiu~O_TRACE_DATA19  = tpiu_TRACE_DATA_bus[19];
assign \tpiu~O_TRACE_DATA20  = tpiu_TRACE_DATA_bus[20];
assign \tpiu~O_TRACE_DATA21  = tpiu_TRACE_DATA_bus[21];
assign \tpiu~O_TRACE_DATA22  = tpiu_TRACE_DATA_bus[22];
assign \tpiu~O_TRACE_DATA23  = tpiu_TRACE_DATA_bus[23];
assign \tpiu~O_TRACE_DATA24  = tpiu_TRACE_DATA_bus[24];
assign \tpiu~O_TRACE_DATA25  = tpiu_TRACE_DATA_bus[25];
assign \tpiu~O_TRACE_DATA26  = tpiu_TRACE_DATA_bus[26];
assign \tpiu~O_TRACE_DATA27  = tpiu_TRACE_DATA_bus[27];
assign \tpiu~O_TRACE_DATA28  = tpiu_TRACE_DATA_bus[28];
assign \tpiu~O_TRACE_DATA29  = tpiu_TRACE_DATA_bus[29];
assign \tpiu~O_TRACE_DATA30  = tpiu_TRACE_DATA_bus[30];
assign \tpiu~O_TRACE_DATA31  = tpiu_TRACE_DATA_bus[31];

assign \h2f_ARADDR[0]  = hps2fpga_ARADDR_bus[0];
assign \h2f_ARADDR[1]  = hps2fpga_ARADDR_bus[1];
assign \h2f_ARADDR[2]  = hps2fpga_ARADDR_bus[2];
assign \h2f_ARADDR[3]  = hps2fpga_ARADDR_bus[3];
assign \h2f_ARADDR[4]  = hps2fpga_ARADDR_bus[4];
assign \h2f_ARADDR[5]  = hps2fpga_ARADDR_bus[5];
assign \h2f_ARADDR[6]  = hps2fpga_ARADDR_bus[6];
assign \h2f_ARADDR[7]  = hps2fpga_ARADDR_bus[7];
assign \h2f_ARADDR[8]  = hps2fpga_ARADDR_bus[8];
assign \h2f_ARADDR[9]  = hps2fpga_ARADDR_bus[9];
assign \h2f_ARADDR[10]  = hps2fpga_ARADDR_bus[10];
assign \h2f_ARADDR[11]  = hps2fpga_ARADDR_bus[11];
assign \h2f_ARADDR[12]  = hps2fpga_ARADDR_bus[12];
assign \h2f_ARADDR[13]  = hps2fpga_ARADDR_bus[13];
assign \h2f_ARADDR[14]  = hps2fpga_ARADDR_bus[14];
assign \h2f_ARADDR[15]  = hps2fpga_ARADDR_bus[15];
assign \h2f_ARADDR[16]  = hps2fpga_ARADDR_bus[16];
assign \h2f_ARADDR[17]  = hps2fpga_ARADDR_bus[17];
assign \h2f_ARADDR[18]  = hps2fpga_ARADDR_bus[18];
assign \h2f_ARADDR[19]  = hps2fpga_ARADDR_bus[19];
assign \h2f_ARADDR[20]  = hps2fpga_ARADDR_bus[20];
assign \h2f_ARADDR[21]  = hps2fpga_ARADDR_bus[21];
assign \h2f_ARADDR[22]  = hps2fpga_ARADDR_bus[22];
assign \h2f_ARADDR[23]  = hps2fpga_ARADDR_bus[23];
assign \h2f_ARADDR[24]  = hps2fpga_ARADDR_bus[24];
assign \h2f_ARADDR[25]  = hps2fpga_ARADDR_bus[25];
assign \h2f_ARADDR[26]  = hps2fpga_ARADDR_bus[26];
assign \h2f_ARADDR[27]  = hps2fpga_ARADDR_bus[27];
assign \h2f_ARADDR[28]  = hps2fpga_ARADDR_bus[28];
assign \h2f_ARADDR[29]  = hps2fpga_ARADDR_bus[29];

assign h2f_lw_ARADDR[0] = hps2fpga_light_weight_ARADDR_bus[0];
assign h2f_lw_ARADDR[1] = hps2fpga_light_weight_ARADDR_bus[1];
assign h2f_lw_ARADDR[2] = hps2fpga_light_weight_ARADDR_bus[2];
assign h2f_lw_ARADDR[3] = hps2fpga_light_weight_ARADDR_bus[3];
assign h2f_lw_ARADDR[4] = hps2fpga_light_weight_ARADDR_bus[4];
assign h2f_lw_ARADDR[5] = hps2fpga_light_weight_ARADDR_bus[5];
assign h2f_lw_ARADDR[6] = hps2fpga_light_weight_ARADDR_bus[6];
assign h2f_lw_ARADDR[7] = hps2fpga_light_weight_ARADDR_bus[7];
assign h2f_lw_ARADDR[8] = hps2fpga_light_weight_ARADDR_bus[8];
assign h2f_lw_ARADDR[9] = hps2fpga_light_weight_ARADDR_bus[9];
assign h2f_lw_ARADDR[10] = hps2fpga_light_weight_ARADDR_bus[10];
assign h2f_lw_ARADDR[11] = hps2fpga_light_weight_ARADDR_bus[11];
assign h2f_lw_ARADDR[12] = hps2fpga_light_weight_ARADDR_bus[12];
assign h2f_lw_ARADDR[13] = hps2fpga_light_weight_ARADDR_bus[13];
assign h2f_lw_ARADDR[14] = hps2fpga_light_weight_ARADDR_bus[14];
assign h2f_lw_ARADDR[15] = hps2fpga_light_weight_ARADDR_bus[15];
assign h2f_lw_ARADDR[16] = hps2fpga_light_weight_ARADDR_bus[16];
assign h2f_lw_ARADDR[17] = hps2fpga_light_weight_ARADDR_bus[17];
assign h2f_lw_ARADDR[18] = hps2fpga_light_weight_ARADDR_bus[18];
assign \h2f_lw_ARADDR[19]  = hps2fpga_light_weight_ARADDR_bus[19];
assign \h2f_lw_ARADDR[20]  = hps2fpga_light_weight_ARADDR_bus[20];

assign h2f_lw_ARBURST[0] = hps2fpga_light_weight_ARBURST_bus[0];
assign h2f_lw_ARBURST[1] = hps2fpga_light_weight_ARBURST_bus[1];

assign h2f_lw_ARID[0] = hps2fpga_light_weight_ARID_bus[0];
assign h2f_lw_ARID[1] = hps2fpga_light_weight_ARID_bus[1];
assign h2f_lw_ARID[2] = hps2fpga_light_weight_ARID_bus[2];
assign h2f_lw_ARID[3] = hps2fpga_light_weight_ARID_bus[3];
assign h2f_lw_ARID[4] = hps2fpga_light_weight_ARID_bus[4];
assign h2f_lw_ARID[5] = hps2fpga_light_weight_ARID_bus[5];
assign h2f_lw_ARID[6] = hps2fpga_light_weight_ARID_bus[6];
assign h2f_lw_ARID[7] = hps2fpga_light_weight_ARID_bus[7];
assign h2f_lw_ARID[8] = hps2fpga_light_weight_ARID_bus[8];
assign h2f_lw_ARID[9] = hps2fpga_light_weight_ARID_bus[9];
assign h2f_lw_ARID[10] = hps2fpga_light_weight_ARID_bus[10];
assign h2f_lw_ARID[11] = hps2fpga_light_weight_ARID_bus[11];

assign h2f_lw_ARLEN[0] = hps2fpga_light_weight_ARLEN_bus[0];
assign h2f_lw_ARLEN[1] = hps2fpga_light_weight_ARLEN_bus[1];
assign h2f_lw_ARLEN[2] = hps2fpga_light_weight_ARLEN_bus[2];
assign h2f_lw_ARLEN[3] = hps2fpga_light_weight_ARLEN_bus[3];

assign h2f_lw_ARSIZE[0] = hps2fpga_light_weight_ARSIZE_bus[0];
assign h2f_lw_ARSIZE[1] = hps2fpga_light_weight_ARSIZE_bus[1];
assign h2f_lw_ARSIZE[2] = hps2fpga_light_weight_ARSIZE_bus[2];

assign h2f_lw_AWADDR[0] = hps2fpga_light_weight_AWADDR_bus[0];
assign h2f_lw_AWADDR[1] = hps2fpga_light_weight_AWADDR_bus[1];
assign h2f_lw_AWADDR[2] = hps2fpga_light_weight_AWADDR_bus[2];
assign h2f_lw_AWADDR[3] = hps2fpga_light_weight_AWADDR_bus[3];
assign h2f_lw_AWADDR[4] = hps2fpga_light_weight_AWADDR_bus[4];
assign h2f_lw_AWADDR[5] = hps2fpga_light_weight_AWADDR_bus[5];
assign h2f_lw_AWADDR[6] = hps2fpga_light_weight_AWADDR_bus[6];
assign h2f_lw_AWADDR[7] = hps2fpga_light_weight_AWADDR_bus[7];
assign h2f_lw_AWADDR[8] = hps2fpga_light_weight_AWADDR_bus[8];
assign h2f_lw_AWADDR[9] = hps2fpga_light_weight_AWADDR_bus[9];
assign h2f_lw_AWADDR[10] = hps2fpga_light_weight_AWADDR_bus[10];
assign h2f_lw_AWADDR[11] = hps2fpga_light_weight_AWADDR_bus[11];
assign h2f_lw_AWADDR[12] = hps2fpga_light_weight_AWADDR_bus[12];
assign h2f_lw_AWADDR[13] = hps2fpga_light_weight_AWADDR_bus[13];
assign h2f_lw_AWADDR[14] = hps2fpga_light_weight_AWADDR_bus[14];
assign h2f_lw_AWADDR[15] = hps2fpga_light_weight_AWADDR_bus[15];
assign h2f_lw_AWADDR[16] = hps2fpga_light_weight_AWADDR_bus[16];
assign h2f_lw_AWADDR[17] = hps2fpga_light_weight_AWADDR_bus[17];
assign h2f_lw_AWADDR[18] = hps2fpga_light_weight_AWADDR_bus[18];

assign h2f_lw_AWBURST[0] = hps2fpga_light_weight_AWBURST_bus[0];
assign h2f_lw_AWBURST[1] = hps2fpga_light_weight_AWBURST_bus[1];

assign h2f_lw_AWID[0] = hps2fpga_light_weight_AWID_bus[0];
assign h2f_lw_AWID[1] = hps2fpga_light_weight_AWID_bus[1];
assign h2f_lw_AWID[2] = hps2fpga_light_weight_AWID_bus[2];
assign h2f_lw_AWID[3] = hps2fpga_light_weight_AWID_bus[3];
assign h2f_lw_AWID[4] = hps2fpga_light_weight_AWID_bus[4];
assign h2f_lw_AWID[5] = hps2fpga_light_weight_AWID_bus[5];
assign h2f_lw_AWID[6] = hps2fpga_light_weight_AWID_bus[6];
assign h2f_lw_AWID[7] = hps2fpga_light_weight_AWID_bus[7];
assign h2f_lw_AWID[8] = hps2fpga_light_weight_AWID_bus[8];
assign h2f_lw_AWID[9] = hps2fpga_light_weight_AWID_bus[9];
assign h2f_lw_AWID[10] = hps2fpga_light_weight_AWID_bus[10];
assign h2f_lw_AWID[11] = hps2fpga_light_weight_AWID_bus[11];

assign h2f_lw_AWLEN[0] = hps2fpga_light_weight_AWLEN_bus[0];
assign h2f_lw_AWLEN[1] = hps2fpga_light_weight_AWLEN_bus[1];
assign h2f_lw_AWLEN[2] = hps2fpga_light_weight_AWLEN_bus[2];
assign h2f_lw_AWLEN[3] = hps2fpga_light_weight_AWLEN_bus[3];

assign h2f_lw_AWSIZE[0] = hps2fpga_light_weight_AWSIZE_bus[0];
assign h2f_lw_AWSIZE[1] = hps2fpga_light_weight_AWSIZE_bus[1];
assign h2f_lw_AWSIZE[2] = hps2fpga_light_weight_AWSIZE_bus[2];

assign h2f_lw_WDATA[0] = hps2fpga_light_weight_WDATA_bus[0];
assign h2f_lw_WDATA[1] = hps2fpga_light_weight_WDATA_bus[1];
assign h2f_lw_WDATA[2] = hps2fpga_light_weight_WDATA_bus[2];
assign h2f_lw_WDATA[3] = hps2fpga_light_weight_WDATA_bus[3];
assign h2f_lw_WDATA[4] = hps2fpga_light_weight_WDATA_bus[4];
assign h2f_lw_WDATA[5] = hps2fpga_light_weight_WDATA_bus[5];
assign h2f_lw_WDATA[6] = hps2fpga_light_weight_WDATA_bus[6];
assign h2f_lw_WDATA[7] = hps2fpga_light_weight_WDATA_bus[7];
assign h2f_lw_WDATA[8] = hps2fpga_light_weight_WDATA_bus[8];
assign h2f_lw_WDATA[9] = hps2fpga_light_weight_WDATA_bus[9];
assign h2f_lw_WDATA[10] = hps2fpga_light_weight_WDATA_bus[10];
assign h2f_lw_WDATA[11] = hps2fpga_light_weight_WDATA_bus[11];
assign h2f_lw_WDATA[12] = hps2fpga_light_weight_WDATA_bus[12];
assign h2f_lw_WDATA[13] = hps2fpga_light_weight_WDATA_bus[13];
assign h2f_lw_WDATA[14] = hps2fpga_light_weight_WDATA_bus[14];
assign h2f_lw_WDATA[15] = hps2fpga_light_weight_WDATA_bus[15];
assign h2f_lw_WDATA[16] = hps2fpga_light_weight_WDATA_bus[16];
assign h2f_lw_WDATA[17] = hps2fpga_light_weight_WDATA_bus[17];
assign h2f_lw_WDATA[18] = hps2fpga_light_weight_WDATA_bus[18];
assign h2f_lw_WDATA[19] = hps2fpga_light_weight_WDATA_bus[19];
assign h2f_lw_WDATA[20] = hps2fpga_light_weight_WDATA_bus[20];
assign h2f_lw_WDATA[21] = hps2fpga_light_weight_WDATA_bus[21];
assign h2f_lw_WDATA[22] = hps2fpga_light_weight_WDATA_bus[22];
assign h2f_lw_WDATA[23] = hps2fpga_light_weight_WDATA_bus[23];
assign h2f_lw_WDATA[24] = hps2fpga_light_weight_WDATA_bus[24];
assign h2f_lw_WDATA[25] = hps2fpga_light_weight_WDATA_bus[25];
assign h2f_lw_WDATA[26] = hps2fpga_light_weight_WDATA_bus[26];
assign h2f_lw_WDATA[27] = hps2fpga_light_weight_WDATA_bus[27];
assign h2f_lw_WDATA[28] = hps2fpga_light_weight_WDATA_bus[28];
assign h2f_lw_WDATA[29] = hps2fpga_light_weight_WDATA_bus[29];
assign h2f_lw_WDATA[30] = hps2fpga_light_weight_WDATA_bus[30];
assign h2f_lw_WDATA[31] = hps2fpga_light_weight_WDATA_bus[31];

assign h2f_lw_WSTRB[0] = hps2fpga_light_weight_WSTRB_bus[0];
assign h2f_lw_WSTRB[1] = hps2fpga_light_weight_WSTRB_bus[1];
assign h2f_lw_WSTRB[2] = hps2fpga_light_weight_WSTRB_bus[2];
assign h2f_lw_WSTRB[3] = hps2fpga_light_weight_WSTRB_bus[3];

assign \f2sdram~O_BONDING_OUT_10  = f2sdram_BONDING_OUT_1_bus[0];
assign \f2sdram~O_BONDING_OUT_11  = f2sdram_BONDING_OUT_1_bus[1];
assign \f2sdram~O_BONDING_OUT_12  = f2sdram_BONDING_OUT_1_bus[2];
assign \f2sdram~O_BONDING_OUT_13  = f2sdram_BONDING_OUT_1_bus[3];

assign f2h_sdram0_READDATA[0] = f2sdram_RD_DATA_0_bus[0];
assign f2h_sdram0_READDATA[1] = f2sdram_RD_DATA_0_bus[1];
assign f2h_sdram0_READDATA[2] = f2sdram_RD_DATA_0_bus[2];
assign f2h_sdram0_READDATA[3] = f2sdram_RD_DATA_0_bus[3];
assign f2h_sdram0_READDATA[4] = f2sdram_RD_DATA_0_bus[4];
assign f2h_sdram0_READDATA[5] = f2sdram_RD_DATA_0_bus[5];
assign f2h_sdram0_READDATA[6] = f2sdram_RD_DATA_0_bus[6];
assign f2h_sdram0_READDATA[7] = f2sdram_RD_DATA_0_bus[7];
assign f2h_sdram0_READDATA[8] = f2sdram_RD_DATA_0_bus[8];
assign f2h_sdram0_READDATA[9] = f2sdram_RD_DATA_0_bus[9];
assign f2h_sdram0_READDATA[10] = f2sdram_RD_DATA_0_bus[10];
assign f2h_sdram0_READDATA[11] = f2sdram_RD_DATA_0_bus[11];
assign f2h_sdram0_READDATA[12] = f2sdram_RD_DATA_0_bus[12];
assign f2h_sdram0_READDATA[13] = f2sdram_RD_DATA_0_bus[13];
assign f2h_sdram0_READDATA[14] = f2sdram_RD_DATA_0_bus[14];
assign f2h_sdram0_READDATA[15] = f2sdram_RD_DATA_0_bus[15];
assign f2h_sdram0_READDATA[16] = f2sdram_RD_DATA_0_bus[16];
assign f2h_sdram0_READDATA[17] = f2sdram_RD_DATA_0_bus[17];
assign f2h_sdram0_READDATA[18] = f2sdram_RD_DATA_0_bus[18];
assign f2h_sdram0_READDATA[19] = f2sdram_RD_DATA_0_bus[19];
assign f2h_sdram0_READDATA[20] = f2sdram_RD_DATA_0_bus[20];
assign f2h_sdram0_READDATA[21] = f2sdram_RD_DATA_0_bus[21];
assign f2h_sdram0_READDATA[22] = f2sdram_RD_DATA_0_bus[22];
assign f2h_sdram0_READDATA[23] = f2sdram_RD_DATA_0_bus[23];
assign f2h_sdram0_READDATA[24] = f2sdram_RD_DATA_0_bus[24];
assign f2h_sdram0_READDATA[25] = f2sdram_RD_DATA_0_bus[25];
assign f2h_sdram0_READDATA[26] = f2sdram_RD_DATA_0_bus[26];
assign f2h_sdram0_READDATA[27] = f2sdram_RD_DATA_0_bus[27];
assign f2h_sdram0_READDATA[28] = f2sdram_RD_DATA_0_bus[28];
assign f2h_sdram0_READDATA[29] = f2sdram_RD_DATA_0_bus[29];
assign f2h_sdram0_READDATA[30] = f2sdram_RD_DATA_0_bus[30];
assign f2h_sdram0_READDATA[31] = f2sdram_RD_DATA_0_bus[31];
assign f2h_sdram0_READDATA[32] = f2sdram_RD_DATA_0_bus[32];
assign f2h_sdram0_READDATA[33] = f2sdram_RD_DATA_0_bus[33];
assign f2h_sdram0_READDATA[34] = f2sdram_RD_DATA_0_bus[34];
assign f2h_sdram0_READDATA[35] = f2sdram_RD_DATA_0_bus[35];
assign f2h_sdram0_READDATA[36] = f2sdram_RD_DATA_0_bus[36];
assign f2h_sdram0_READDATA[37] = f2sdram_RD_DATA_0_bus[37];
assign f2h_sdram0_READDATA[38] = f2sdram_RD_DATA_0_bus[38];
assign f2h_sdram0_READDATA[39] = f2sdram_RD_DATA_0_bus[39];
assign f2h_sdram0_READDATA[40] = f2sdram_RD_DATA_0_bus[40];
assign f2h_sdram0_READDATA[41] = f2sdram_RD_DATA_0_bus[41];
assign f2h_sdram0_READDATA[42] = f2sdram_RD_DATA_0_bus[42];
assign f2h_sdram0_READDATA[43] = f2sdram_RD_DATA_0_bus[43];
assign f2h_sdram0_READDATA[44] = f2sdram_RD_DATA_0_bus[44];
assign f2h_sdram0_READDATA[45] = f2sdram_RD_DATA_0_bus[45];
assign f2h_sdram0_READDATA[46] = f2sdram_RD_DATA_0_bus[46];
assign f2h_sdram0_READDATA[47] = f2sdram_RD_DATA_0_bus[47];
assign f2h_sdram0_READDATA[48] = f2sdram_RD_DATA_0_bus[48];
assign f2h_sdram0_READDATA[49] = f2sdram_RD_DATA_0_bus[49];
assign f2h_sdram0_READDATA[50] = f2sdram_RD_DATA_0_bus[50];
assign f2h_sdram0_READDATA[51] = f2sdram_RD_DATA_0_bus[51];
assign f2h_sdram0_READDATA[52] = f2sdram_RD_DATA_0_bus[52];
assign f2h_sdram0_READDATA[53] = f2sdram_RD_DATA_0_bus[53];
assign f2h_sdram0_READDATA[54] = f2sdram_RD_DATA_0_bus[54];
assign f2h_sdram0_READDATA[55] = f2sdram_RD_DATA_0_bus[55];
assign f2h_sdram0_READDATA[56] = f2sdram_RD_DATA_0_bus[56];
assign f2h_sdram0_READDATA[57] = f2sdram_RD_DATA_0_bus[57];
assign f2h_sdram0_READDATA[58] = f2sdram_RD_DATA_0_bus[58];
assign f2h_sdram0_READDATA[59] = f2sdram_RD_DATA_0_bus[59];
assign f2h_sdram0_READDATA[60] = f2sdram_RD_DATA_0_bus[60];
assign f2h_sdram0_READDATA[61] = f2sdram_RD_DATA_0_bus[61];
assign f2h_sdram0_READDATA[62] = f2sdram_RD_DATA_0_bus[62];
assign f2h_sdram0_READDATA[63] = f2sdram_RD_DATA_0_bus[63];

assign f2h_sdram0_READDATA[64] = f2sdram_RD_DATA_1_bus[0];
assign f2h_sdram0_READDATA[65] = f2sdram_RD_DATA_1_bus[1];
assign f2h_sdram0_READDATA[66] = f2sdram_RD_DATA_1_bus[2];
assign f2h_sdram0_READDATA[67] = f2sdram_RD_DATA_1_bus[3];
assign f2h_sdram0_READDATA[68] = f2sdram_RD_DATA_1_bus[4];
assign f2h_sdram0_READDATA[69] = f2sdram_RD_DATA_1_bus[5];
assign f2h_sdram0_READDATA[70] = f2sdram_RD_DATA_1_bus[6];
assign f2h_sdram0_READDATA[71] = f2sdram_RD_DATA_1_bus[7];
assign f2h_sdram0_READDATA[72] = f2sdram_RD_DATA_1_bus[8];
assign f2h_sdram0_READDATA[73] = f2sdram_RD_DATA_1_bus[9];
assign f2h_sdram0_READDATA[74] = f2sdram_RD_DATA_1_bus[10];
assign f2h_sdram0_READDATA[75] = f2sdram_RD_DATA_1_bus[11];
assign f2h_sdram0_READDATA[76] = f2sdram_RD_DATA_1_bus[12];
assign f2h_sdram0_READDATA[77] = f2sdram_RD_DATA_1_bus[13];
assign f2h_sdram0_READDATA[78] = f2sdram_RD_DATA_1_bus[14];
assign f2h_sdram0_READDATA[79] = f2sdram_RD_DATA_1_bus[15];
assign f2h_sdram0_READDATA[80] = f2sdram_RD_DATA_1_bus[16];
assign f2h_sdram0_READDATA[81] = f2sdram_RD_DATA_1_bus[17];
assign f2h_sdram0_READDATA[82] = f2sdram_RD_DATA_1_bus[18];
assign f2h_sdram0_READDATA[83] = f2sdram_RD_DATA_1_bus[19];
assign f2h_sdram0_READDATA[84] = f2sdram_RD_DATA_1_bus[20];
assign f2h_sdram0_READDATA[85] = f2sdram_RD_DATA_1_bus[21];
assign f2h_sdram0_READDATA[86] = f2sdram_RD_DATA_1_bus[22];
assign f2h_sdram0_READDATA[87] = f2sdram_RD_DATA_1_bus[23];
assign f2h_sdram0_READDATA[88] = f2sdram_RD_DATA_1_bus[24];
assign f2h_sdram0_READDATA[89] = f2sdram_RD_DATA_1_bus[25];
assign f2h_sdram0_READDATA[90] = f2sdram_RD_DATA_1_bus[26];
assign f2h_sdram0_READDATA[91] = f2sdram_RD_DATA_1_bus[27];
assign f2h_sdram0_READDATA[92] = f2sdram_RD_DATA_1_bus[28];
assign f2h_sdram0_READDATA[93] = f2sdram_RD_DATA_1_bus[29];
assign f2h_sdram0_READDATA[94] = f2sdram_RD_DATA_1_bus[30];
assign f2h_sdram0_READDATA[95] = f2sdram_RD_DATA_1_bus[31];
assign f2h_sdram0_READDATA[96] = f2sdram_RD_DATA_1_bus[32];
assign f2h_sdram0_READDATA[97] = f2sdram_RD_DATA_1_bus[33];
assign f2h_sdram0_READDATA[98] = f2sdram_RD_DATA_1_bus[34];
assign f2h_sdram0_READDATA[99] = f2sdram_RD_DATA_1_bus[35];
assign f2h_sdram0_READDATA[100] = f2sdram_RD_DATA_1_bus[36];
assign f2h_sdram0_READDATA[101] = f2sdram_RD_DATA_1_bus[37];
assign f2h_sdram0_READDATA[102] = f2sdram_RD_DATA_1_bus[38];
assign f2h_sdram0_READDATA[103] = f2sdram_RD_DATA_1_bus[39];
assign f2h_sdram0_READDATA[104] = f2sdram_RD_DATA_1_bus[40];
assign f2h_sdram0_READDATA[105] = f2sdram_RD_DATA_1_bus[41];
assign f2h_sdram0_READDATA[106] = f2sdram_RD_DATA_1_bus[42];
assign f2h_sdram0_READDATA[107] = f2sdram_RD_DATA_1_bus[43];
assign f2h_sdram0_READDATA[108] = f2sdram_RD_DATA_1_bus[44];
assign f2h_sdram0_READDATA[109] = f2sdram_RD_DATA_1_bus[45];
assign f2h_sdram0_READDATA[110] = f2sdram_RD_DATA_1_bus[46];
assign f2h_sdram0_READDATA[111] = f2sdram_RD_DATA_1_bus[47];
assign f2h_sdram0_READDATA[112] = f2sdram_RD_DATA_1_bus[48];
assign f2h_sdram0_READDATA[113] = f2sdram_RD_DATA_1_bus[49];
assign f2h_sdram0_READDATA[114] = f2sdram_RD_DATA_1_bus[50];
assign f2h_sdram0_READDATA[115] = f2sdram_RD_DATA_1_bus[51];
assign f2h_sdram0_READDATA[116] = f2sdram_RD_DATA_1_bus[52];
assign f2h_sdram0_READDATA[117] = f2sdram_RD_DATA_1_bus[53];
assign f2h_sdram0_READDATA[118] = f2sdram_RD_DATA_1_bus[54];
assign f2h_sdram0_READDATA[119] = f2sdram_RD_DATA_1_bus[55];
assign f2h_sdram0_READDATA[120] = f2sdram_RD_DATA_1_bus[56];
assign f2h_sdram0_READDATA[121] = f2sdram_RD_DATA_1_bus[57];
assign f2h_sdram0_READDATA[122] = f2sdram_RD_DATA_1_bus[58];
assign f2h_sdram0_READDATA[123] = f2sdram_RD_DATA_1_bus[59];
assign f2h_sdram0_READDATA[124] = f2sdram_RD_DATA_1_bus[60];
assign f2h_sdram0_READDATA[125] = f2sdram_RD_DATA_1_bus[61];
assign f2h_sdram0_READDATA[126] = f2sdram_RD_DATA_1_bus[62];
assign f2h_sdram0_READDATA[127] = f2sdram_RD_DATA_1_bus[63];

assign f2h_sdram0_READDATA[128] = f2sdram_RD_DATA_2_bus[0];
assign f2h_sdram0_READDATA[129] = f2sdram_RD_DATA_2_bus[1];
assign f2h_sdram0_READDATA[130] = f2sdram_RD_DATA_2_bus[2];
assign f2h_sdram0_READDATA[131] = f2sdram_RD_DATA_2_bus[3];
assign f2h_sdram0_READDATA[132] = f2sdram_RD_DATA_2_bus[4];
assign f2h_sdram0_READDATA[133] = f2sdram_RD_DATA_2_bus[5];
assign f2h_sdram0_READDATA[134] = f2sdram_RD_DATA_2_bus[6];
assign f2h_sdram0_READDATA[135] = f2sdram_RD_DATA_2_bus[7];
assign f2h_sdram0_READDATA[136] = f2sdram_RD_DATA_2_bus[8];
assign f2h_sdram0_READDATA[137] = f2sdram_RD_DATA_2_bus[9];
assign f2h_sdram0_READDATA[138] = f2sdram_RD_DATA_2_bus[10];
assign f2h_sdram0_READDATA[139] = f2sdram_RD_DATA_2_bus[11];
assign f2h_sdram0_READDATA[140] = f2sdram_RD_DATA_2_bus[12];
assign f2h_sdram0_READDATA[141] = f2sdram_RD_DATA_2_bus[13];
assign f2h_sdram0_READDATA[142] = f2sdram_RD_DATA_2_bus[14];
assign f2h_sdram0_READDATA[143] = f2sdram_RD_DATA_2_bus[15];
assign f2h_sdram0_READDATA[144] = f2sdram_RD_DATA_2_bus[16];
assign f2h_sdram0_READDATA[145] = f2sdram_RD_DATA_2_bus[17];
assign f2h_sdram0_READDATA[146] = f2sdram_RD_DATA_2_bus[18];
assign f2h_sdram0_READDATA[147] = f2sdram_RD_DATA_2_bus[19];
assign f2h_sdram0_READDATA[148] = f2sdram_RD_DATA_2_bus[20];
assign f2h_sdram0_READDATA[149] = f2sdram_RD_DATA_2_bus[21];
assign f2h_sdram0_READDATA[150] = f2sdram_RD_DATA_2_bus[22];
assign f2h_sdram0_READDATA[151] = f2sdram_RD_DATA_2_bus[23];
assign f2h_sdram0_READDATA[152] = f2sdram_RD_DATA_2_bus[24];
assign f2h_sdram0_READDATA[153] = f2sdram_RD_DATA_2_bus[25];
assign f2h_sdram0_READDATA[154] = f2sdram_RD_DATA_2_bus[26];
assign f2h_sdram0_READDATA[155] = f2sdram_RD_DATA_2_bus[27];
assign f2h_sdram0_READDATA[156] = f2sdram_RD_DATA_2_bus[28];
assign f2h_sdram0_READDATA[157] = f2sdram_RD_DATA_2_bus[29];
assign f2h_sdram0_READDATA[158] = f2sdram_RD_DATA_2_bus[30];
assign f2h_sdram0_READDATA[159] = f2sdram_RD_DATA_2_bus[31];
assign f2h_sdram0_READDATA[160] = f2sdram_RD_DATA_2_bus[32];
assign f2h_sdram0_READDATA[161] = f2sdram_RD_DATA_2_bus[33];
assign f2h_sdram0_READDATA[162] = f2sdram_RD_DATA_2_bus[34];
assign f2h_sdram0_READDATA[163] = f2sdram_RD_DATA_2_bus[35];
assign f2h_sdram0_READDATA[164] = f2sdram_RD_DATA_2_bus[36];
assign f2h_sdram0_READDATA[165] = f2sdram_RD_DATA_2_bus[37];
assign f2h_sdram0_READDATA[166] = f2sdram_RD_DATA_2_bus[38];
assign f2h_sdram0_READDATA[167] = f2sdram_RD_DATA_2_bus[39];
assign f2h_sdram0_READDATA[168] = f2sdram_RD_DATA_2_bus[40];
assign f2h_sdram0_READDATA[169] = f2sdram_RD_DATA_2_bus[41];
assign f2h_sdram0_READDATA[170] = f2sdram_RD_DATA_2_bus[42];
assign f2h_sdram0_READDATA[171] = f2sdram_RD_DATA_2_bus[43];
assign f2h_sdram0_READDATA[172] = f2sdram_RD_DATA_2_bus[44];
assign f2h_sdram0_READDATA[173] = f2sdram_RD_DATA_2_bus[45];
assign f2h_sdram0_READDATA[174] = f2sdram_RD_DATA_2_bus[46];
assign f2h_sdram0_READDATA[175] = f2sdram_RD_DATA_2_bus[47];
assign f2h_sdram0_READDATA[176] = f2sdram_RD_DATA_2_bus[48];
assign f2h_sdram0_READDATA[177] = f2sdram_RD_DATA_2_bus[49];
assign f2h_sdram0_READDATA[178] = f2sdram_RD_DATA_2_bus[50];
assign f2h_sdram0_READDATA[179] = f2sdram_RD_DATA_2_bus[51];
assign f2h_sdram0_READDATA[180] = f2sdram_RD_DATA_2_bus[52];
assign f2h_sdram0_READDATA[181] = f2sdram_RD_DATA_2_bus[53];
assign f2h_sdram0_READDATA[182] = f2sdram_RD_DATA_2_bus[54];
assign f2h_sdram0_READDATA[183] = f2sdram_RD_DATA_2_bus[55];
assign f2h_sdram0_READDATA[184] = f2sdram_RD_DATA_2_bus[56];
assign f2h_sdram0_READDATA[185] = f2sdram_RD_DATA_2_bus[57];
assign f2h_sdram0_READDATA[186] = f2sdram_RD_DATA_2_bus[58];
assign f2h_sdram0_READDATA[187] = f2sdram_RD_DATA_2_bus[59];
assign f2h_sdram0_READDATA[188] = f2sdram_RD_DATA_2_bus[60];
assign f2h_sdram0_READDATA[189] = f2sdram_RD_DATA_2_bus[61];
assign f2h_sdram0_READDATA[190] = f2sdram_RD_DATA_2_bus[62];
assign f2h_sdram0_READDATA[191] = f2sdram_RD_DATA_2_bus[63];

assign f2h_sdram0_READDATA[192] = f2sdram_RD_DATA_3_bus[0];
assign f2h_sdram0_READDATA[193] = f2sdram_RD_DATA_3_bus[1];
assign f2h_sdram0_READDATA[194] = f2sdram_RD_DATA_3_bus[2];
assign f2h_sdram0_READDATA[195] = f2sdram_RD_DATA_3_bus[3];
assign f2h_sdram0_READDATA[196] = f2sdram_RD_DATA_3_bus[4];
assign f2h_sdram0_READDATA[197] = f2sdram_RD_DATA_3_bus[5];
assign f2h_sdram0_READDATA[198] = f2sdram_RD_DATA_3_bus[6];
assign f2h_sdram0_READDATA[199] = f2sdram_RD_DATA_3_bus[7];
assign f2h_sdram0_READDATA[200] = f2sdram_RD_DATA_3_bus[8];
assign f2h_sdram0_READDATA[201] = f2sdram_RD_DATA_3_bus[9];
assign f2h_sdram0_READDATA[202] = f2sdram_RD_DATA_3_bus[10];
assign f2h_sdram0_READDATA[203] = f2sdram_RD_DATA_3_bus[11];
assign f2h_sdram0_READDATA[204] = f2sdram_RD_DATA_3_bus[12];
assign f2h_sdram0_READDATA[205] = f2sdram_RD_DATA_3_bus[13];
assign f2h_sdram0_READDATA[206] = f2sdram_RD_DATA_3_bus[14];
assign f2h_sdram0_READDATA[207] = f2sdram_RD_DATA_3_bus[15];
assign f2h_sdram0_READDATA[208] = f2sdram_RD_DATA_3_bus[16];
assign f2h_sdram0_READDATA[209] = f2sdram_RD_DATA_3_bus[17];
assign f2h_sdram0_READDATA[210] = f2sdram_RD_DATA_3_bus[18];
assign f2h_sdram0_READDATA[211] = f2sdram_RD_DATA_3_bus[19];
assign f2h_sdram0_READDATA[212] = f2sdram_RD_DATA_3_bus[20];
assign f2h_sdram0_READDATA[213] = f2sdram_RD_DATA_3_bus[21];
assign f2h_sdram0_READDATA[214] = f2sdram_RD_DATA_3_bus[22];
assign f2h_sdram0_READDATA[215] = f2sdram_RD_DATA_3_bus[23];
assign f2h_sdram0_READDATA[216] = f2sdram_RD_DATA_3_bus[24];
assign f2h_sdram0_READDATA[217] = f2sdram_RD_DATA_3_bus[25];
assign f2h_sdram0_READDATA[218] = f2sdram_RD_DATA_3_bus[26];
assign f2h_sdram0_READDATA[219] = f2sdram_RD_DATA_3_bus[27];
assign f2h_sdram0_READDATA[220] = f2sdram_RD_DATA_3_bus[28];
assign f2h_sdram0_READDATA[221] = f2sdram_RD_DATA_3_bus[29];
assign f2h_sdram0_READDATA[222] = f2sdram_RD_DATA_3_bus[30];
assign f2h_sdram0_READDATA[223] = f2sdram_RD_DATA_3_bus[31];
assign f2h_sdram0_READDATA[224] = f2sdram_RD_DATA_3_bus[32];
assign f2h_sdram0_READDATA[225] = f2sdram_RD_DATA_3_bus[33];
assign f2h_sdram0_READDATA[226] = f2sdram_RD_DATA_3_bus[34];
assign f2h_sdram0_READDATA[227] = f2sdram_RD_DATA_3_bus[35];
assign f2h_sdram0_READDATA[228] = f2sdram_RD_DATA_3_bus[36];
assign f2h_sdram0_READDATA[229] = f2sdram_RD_DATA_3_bus[37];
assign f2h_sdram0_READDATA[230] = f2sdram_RD_DATA_3_bus[38];
assign f2h_sdram0_READDATA[231] = f2sdram_RD_DATA_3_bus[39];
assign f2h_sdram0_READDATA[232] = f2sdram_RD_DATA_3_bus[40];
assign f2h_sdram0_READDATA[233] = f2sdram_RD_DATA_3_bus[41];
assign f2h_sdram0_READDATA[234] = f2sdram_RD_DATA_3_bus[42];
assign f2h_sdram0_READDATA[235] = f2sdram_RD_DATA_3_bus[43];
assign f2h_sdram0_READDATA[236] = f2sdram_RD_DATA_3_bus[44];
assign f2h_sdram0_READDATA[237] = f2sdram_RD_DATA_3_bus[45];
assign f2h_sdram0_READDATA[238] = f2sdram_RD_DATA_3_bus[46];
assign f2h_sdram0_READDATA[239] = f2sdram_RD_DATA_3_bus[47];
assign f2h_sdram0_READDATA[240] = f2sdram_RD_DATA_3_bus[48];
assign f2h_sdram0_READDATA[241] = f2sdram_RD_DATA_3_bus[49];
assign f2h_sdram0_READDATA[242] = f2sdram_RD_DATA_3_bus[50];
assign f2h_sdram0_READDATA[243] = f2sdram_RD_DATA_3_bus[51];
assign f2h_sdram0_READDATA[244] = f2sdram_RD_DATA_3_bus[52];
assign f2h_sdram0_READDATA[245] = f2sdram_RD_DATA_3_bus[53];
assign f2h_sdram0_READDATA[246] = f2sdram_RD_DATA_3_bus[54];
assign f2h_sdram0_READDATA[247] = f2sdram_RD_DATA_3_bus[55];
assign f2h_sdram0_READDATA[248] = f2sdram_RD_DATA_3_bus[56];
assign f2h_sdram0_READDATA[249] = f2sdram_RD_DATA_3_bus[57];
assign f2h_sdram0_READDATA[250] = f2sdram_RD_DATA_3_bus[58];
assign f2h_sdram0_READDATA[251] = f2sdram_RD_DATA_3_bus[59];
assign f2h_sdram0_READDATA[252] = f2sdram_RD_DATA_3_bus[60];
assign f2h_sdram0_READDATA[253] = f2sdram_RD_DATA_3_bus[61];
assign f2h_sdram0_READDATA[254] = f2sdram_RD_DATA_3_bus[62];
assign f2h_sdram0_READDATA[255] = f2sdram_RD_DATA_3_bus[63];

cyclonev_hps_interface_clocks_resets clocks_resets(
	.f2h_cold_rst_req_n(vcc),
	.f2h_dbg_rst_req_n(vcc),
	.f2h_pending_rst_ack(f2h_pending_rst_ack_n[0]),
	.f2h_periph_ref_clk(gnd),
	.f2h_sdram_ref_clk(gnd),
	.f2h_warm_rst_req_n(vcc),
	.ptp_ref_clk(gnd),
	.h2f_cold_rst_n(h2f_cold_rst_n[0]),
	.h2f_pending_rst_req_n(h2f_pending_rst_req_n[0]),
	.h2f_rst_n(h2f_rst_n[0]),
	.h2f_user0_clk(),
	.h2f_user1_clk(),
	.h2f_user2_clk());
defparam clocks_resets.h2f_user0_clk_freq = 100;
defparam clocks_resets.h2f_user1_clk_freq = 100;
defparam clocks_resets.h2f_user2_clk_freq = 100;

cyclonev_hps_interface_hps2fpga_light_weight hps2fpga_light_weight(
	.arready(h2f_lw_ARREADY[0]),
	.awready(h2f_lw_AWREADY[0]),
	.bvalid(h2f_lw_BVALID[0]),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(h2f_lw_RLAST[0]),
	.rvalid(h2f_lw_RVALID[0]),
	.wready(h2f_lw_WREADY[0]),
	.bid({h2f_lw_BID[11],h2f_lw_BID[10],h2f_lw_BID[9],h2f_lw_BID[8],h2f_lw_BID[7],h2f_lw_BID[6],h2f_lw_BID[5],h2f_lw_BID[4],h2f_lw_BID[3],h2f_lw_BID[2],h2f_lw_BID[1],h2f_lw_BID[0]}),
	.bresp({gnd,gnd}),
	.rdata({h2f_lw_RDATA[31],h2f_lw_RDATA[30],h2f_lw_RDATA[29],h2f_lw_RDATA[28],h2f_lw_RDATA[27],h2f_lw_RDATA[26],h2f_lw_RDATA[25],h2f_lw_RDATA[24],h2f_lw_RDATA[23],h2f_lw_RDATA[22],h2f_lw_RDATA[21],h2f_lw_RDATA[20],h2f_lw_RDATA[19],h2f_lw_RDATA[18],h2f_lw_RDATA[17],h2f_lw_RDATA[16],h2f_lw_RDATA[15],h2f_lw_RDATA[14],h2f_lw_RDATA[13],h2f_lw_RDATA[12],h2f_lw_RDATA[11],
h2f_lw_RDATA[10],h2f_lw_RDATA[9],h2f_lw_RDATA[8],h2f_lw_RDATA[7],h2f_lw_RDATA[6],h2f_lw_RDATA[5],h2f_lw_RDATA[4],h2f_lw_RDATA[3],h2f_lw_RDATA[2],h2f_lw_RDATA[1],h2f_lw_RDATA[0]}),
	.rid({h2f_lw_RID[11],h2f_lw_RID[10],h2f_lw_RID[9],h2f_lw_RID[8],h2f_lw_RID[7],h2f_lw_RID[6],h2f_lw_RID[5],h2f_lw_RID[4],h2f_lw_RID[3],h2f_lw_RID[2],h2f_lw_RID[1],h2f_lw_RID[0]}),
	.rresp({gnd,gnd}),
	.arvalid(h2f_lw_ARVALID[0]),
	.awvalid(h2f_lw_AWVALID[0]),
	.bready(h2f_lw_BREADY[0]),
	.rready(h2f_lw_RREADY[0]),
	.wlast(h2f_lw_WLAST[0]),
	.wvalid(h2f_lw_WVALID[0]),
	.araddr(hps2fpga_light_weight_ARADDR_bus),
	.arburst(hps2fpga_light_weight_ARBURST_bus),
	.arcache(),
	.arid(hps2fpga_light_weight_ARID_bus),
	.arlen(hps2fpga_light_weight_ARLEN_bus),
	.arlock(),
	.arprot(),
	.arsize(hps2fpga_light_weight_ARSIZE_bus),
	.awaddr(hps2fpga_light_weight_AWADDR_bus),
	.awburst(hps2fpga_light_weight_AWBURST_bus),
	.awcache(),
	.awid(hps2fpga_light_weight_AWID_bus),
	.awlen(hps2fpga_light_weight_AWLEN_bus),
	.awlock(),
	.awprot(),
	.awsize(hps2fpga_light_weight_AWSIZE_bus),
	.wdata(hps2fpga_light_weight_WDATA_bus),
	.wid(),
	.wstrb(hps2fpga_light_weight_WSTRB_bus));

cyclonev_hps_interface_fpga2sdram f2sdram(
	.cmd_port_clk_0(h2f_lw_axi_clk[0]),
	.cmd_port_clk_1(gnd),
	.cmd_port_clk_2(gnd),
	.cmd_port_clk_3(gnd),
	.cmd_port_clk_4(gnd),
	.cmd_port_clk_5(gnd),
	.cmd_valid_0(\intermediate[12]~combout ),
	.cmd_valid_1(gnd),
	.cmd_valid_2(gnd),
	.cmd_valid_3(gnd),
	.cmd_valid_4(gnd),
	.cmd_valid_5(gnd),
	.rd_clk_0(h2f_lw_axi_clk[0]),
	.rd_clk_1(h2f_lw_axi_clk[0]),
	.rd_clk_2(h2f_lw_axi_clk[0]),
	.rd_clk_3(h2f_lw_axi_clk[0]),
	.rd_ready_0(vcc),
	.rd_ready_1(vcc),
	.rd_ready_2(vcc),
	.rd_ready_3(vcc),
	.wr_clk_0(h2f_lw_axi_clk[0]),
	.wr_clk_1(h2f_lw_axi_clk[0]),
	.wr_clk_2(h2f_lw_axi_clk[0]),
	.wr_clk_3(h2f_lw_axi_clk[0]),
	.wr_valid_0(gnd),
	.wr_valid_1(gnd),
	.wr_valid_2(gnd),
	.wr_valid_3(gnd),
	.wrack_ready_0(vcc),
	.wrack_ready_1(gnd),
	.wrack_ready_2(gnd),
	.wrack_ready_3(gnd),
	.wrack_ready_4(gnd),
	.wrack_ready_5(gnd),
	.cfg_axi_mm_select({gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_rfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_cport_type({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc,vcc}),
	.cfg_cport_wfifo_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_port_width({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,vcc,vcc}),
	.cfg_rfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfg_wfifo_cport_map({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_data_0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_sdram0_BURSTCOUNT[7],f2h_sdram0_BURSTCOUNT[6],f2h_sdram0_BURSTCOUNT[5],f2h_sdram0_BURSTCOUNT[4],f2h_sdram0_BURSTCOUNT[3],f2h_sdram0_BURSTCOUNT[2],f2h_sdram0_BURSTCOUNT[1],f2h_sdram0_BURSTCOUNT[0],gnd,gnd,gnd,gnd,gnd,f2h_sdram0_ADDRESS[26],
f2h_sdram0_ADDRESS[25],f2h_sdram0_ADDRESS[24],f2h_sdram0_ADDRESS[23],f2h_sdram0_ADDRESS[22],f2h_sdram0_ADDRESS[21],f2h_sdram0_ADDRESS[20],f2h_sdram0_ADDRESS[19],f2h_sdram0_ADDRESS[18],f2h_sdram0_ADDRESS[17],f2h_sdram0_ADDRESS[16],f2h_sdram0_ADDRESS[15],f2h_sdram0_ADDRESS[14],f2h_sdram0_ADDRESS[13],f2h_sdram0_ADDRESS[12],
f2h_sdram0_ADDRESS[11],f2h_sdram0_ADDRESS[10],f2h_sdram0_ADDRESS[9],f2h_sdram0_ADDRESS[8],f2h_sdram0_ADDRESS[7],f2h_sdram0_ADDRESS[6],f2h_sdram0_ADDRESS[5],f2h_sdram0_ADDRESS[4],f2h_sdram0_ADDRESS[3],f2h_sdram0_ADDRESS[2],f2h_sdram0_ADDRESS[1],f2h_sdram0_ADDRESS[0],f2h_sdram0_WRITE[0],f2h_sdram0_READ[0]}),
	.cmd_data_1(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_2(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_3(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_4(60'b000000000000000000000000000000000000000000000000000000000000),
	.cmd_data_5(60'b000000000000000000000000000000000000000000000000000000000000),
	.wr_data_0({gnd,gnd,f2h_sdram0_BYTEENABLE[7],f2h_sdram0_BYTEENABLE[6],f2h_sdram0_BYTEENABLE[5],f2h_sdram0_BYTEENABLE[4],f2h_sdram0_BYTEENABLE[3],f2h_sdram0_BYTEENABLE[2],f2h_sdram0_BYTEENABLE[1],f2h_sdram0_BYTEENABLE[0],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_sdram0_WRITEDATA[63],
f2h_sdram0_WRITEDATA[62],f2h_sdram0_WRITEDATA[61],f2h_sdram0_WRITEDATA[60],f2h_sdram0_WRITEDATA[59],f2h_sdram0_WRITEDATA[58],f2h_sdram0_WRITEDATA[57],f2h_sdram0_WRITEDATA[56],f2h_sdram0_WRITEDATA[55],f2h_sdram0_WRITEDATA[54],f2h_sdram0_WRITEDATA[53],f2h_sdram0_WRITEDATA[52],f2h_sdram0_WRITEDATA[51],
f2h_sdram0_WRITEDATA[50],f2h_sdram0_WRITEDATA[49],f2h_sdram0_WRITEDATA[48],f2h_sdram0_WRITEDATA[47],f2h_sdram0_WRITEDATA[46],f2h_sdram0_WRITEDATA[45],f2h_sdram0_WRITEDATA[44],f2h_sdram0_WRITEDATA[43],f2h_sdram0_WRITEDATA[42],f2h_sdram0_WRITEDATA[41],f2h_sdram0_WRITEDATA[40],f2h_sdram0_WRITEDATA[39],
f2h_sdram0_WRITEDATA[38],f2h_sdram0_WRITEDATA[37],f2h_sdram0_WRITEDATA[36],f2h_sdram0_WRITEDATA[35],f2h_sdram0_WRITEDATA[34],f2h_sdram0_WRITEDATA[33],f2h_sdram0_WRITEDATA[32],f2h_sdram0_WRITEDATA[31],f2h_sdram0_WRITEDATA[30],f2h_sdram0_WRITEDATA[29],f2h_sdram0_WRITEDATA[28],f2h_sdram0_WRITEDATA[27],
f2h_sdram0_WRITEDATA[26],f2h_sdram0_WRITEDATA[25],f2h_sdram0_WRITEDATA[24],f2h_sdram0_WRITEDATA[23],f2h_sdram0_WRITEDATA[22],f2h_sdram0_WRITEDATA[21],f2h_sdram0_WRITEDATA[20],f2h_sdram0_WRITEDATA[19],f2h_sdram0_WRITEDATA[18],f2h_sdram0_WRITEDATA[17],f2h_sdram0_WRITEDATA[16],f2h_sdram0_WRITEDATA[15],
f2h_sdram0_WRITEDATA[14],f2h_sdram0_WRITEDATA[13],f2h_sdram0_WRITEDATA[12],f2h_sdram0_WRITEDATA[11],f2h_sdram0_WRITEDATA[10],f2h_sdram0_WRITEDATA[9],f2h_sdram0_WRITEDATA[8],f2h_sdram0_WRITEDATA[7],f2h_sdram0_WRITEDATA[6],f2h_sdram0_WRITEDATA[5],f2h_sdram0_WRITEDATA[4],f2h_sdram0_WRITEDATA[3],
f2h_sdram0_WRITEDATA[2],f2h_sdram0_WRITEDATA[1],f2h_sdram0_WRITEDATA[0]}),
	.wr_data_1({gnd,gnd,f2h_sdram0_BYTEENABLE[15],f2h_sdram0_BYTEENABLE[14],f2h_sdram0_BYTEENABLE[13],f2h_sdram0_BYTEENABLE[12],f2h_sdram0_BYTEENABLE[11],f2h_sdram0_BYTEENABLE[10],f2h_sdram0_BYTEENABLE[9],f2h_sdram0_BYTEENABLE[8],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_sdram0_WRITEDATA[127],
f2h_sdram0_WRITEDATA[126],f2h_sdram0_WRITEDATA[125],f2h_sdram0_WRITEDATA[124],f2h_sdram0_WRITEDATA[123],f2h_sdram0_WRITEDATA[122],f2h_sdram0_WRITEDATA[121],f2h_sdram0_WRITEDATA[120],f2h_sdram0_WRITEDATA[119],f2h_sdram0_WRITEDATA[118],f2h_sdram0_WRITEDATA[117],f2h_sdram0_WRITEDATA[116],f2h_sdram0_WRITEDATA[115],
f2h_sdram0_WRITEDATA[114],f2h_sdram0_WRITEDATA[113],f2h_sdram0_WRITEDATA[112],f2h_sdram0_WRITEDATA[111],f2h_sdram0_WRITEDATA[110],f2h_sdram0_WRITEDATA[109],f2h_sdram0_WRITEDATA[108],f2h_sdram0_WRITEDATA[107],f2h_sdram0_WRITEDATA[106],f2h_sdram0_WRITEDATA[105],f2h_sdram0_WRITEDATA[104],f2h_sdram0_WRITEDATA[103],
f2h_sdram0_WRITEDATA[102],f2h_sdram0_WRITEDATA[101],f2h_sdram0_WRITEDATA[100],f2h_sdram0_WRITEDATA[99],f2h_sdram0_WRITEDATA[98],f2h_sdram0_WRITEDATA[97],f2h_sdram0_WRITEDATA[96],f2h_sdram0_WRITEDATA[95],f2h_sdram0_WRITEDATA[94],f2h_sdram0_WRITEDATA[93],f2h_sdram0_WRITEDATA[92],f2h_sdram0_WRITEDATA[91],
f2h_sdram0_WRITEDATA[90],f2h_sdram0_WRITEDATA[89],f2h_sdram0_WRITEDATA[88],f2h_sdram0_WRITEDATA[87],f2h_sdram0_WRITEDATA[86],f2h_sdram0_WRITEDATA[85],f2h_sdram0_WRITEDATA[84],f2h_sdram0_WRITEDATA[83],f2h_sdram0_WRITEDATA[82],f2h_sdram0_WRITEDATA[81],f2h_sdram0_WRITEDATA[80],f2h_sdram0_WRITEDATA[79],
f2h_sdram0_WRITEDATA[78],f2h_sdram0_WRITEDATA[77],f2h_sdram0_WRITEDATA[76],f2h_sdram0_WRITEDATA[75],f2h_sdram0_WRITEDATA[74],f2h_sdram0_WRITEDATA[73],f2h_sdram0_WRITEDATA[72],f2h_sdram0_WRITEDATA[71],f2h_sdram0_WRITEDATA[70],f2h_sdram0_WRITEDATA[69],f2h_sdram0_WRITEDATA[68],f2h_sdram0_WRITEDATA[67],
f2h_sdram0_WRITEDATA[66],f2h_sdram0_WRITEDATA[65],f2h_sdram0_WRITEDATA[64]}),
	.wr_data_2({gnd,gnd,f2h_sdram0_BYTEENABLE[23],f2h_sdram0_BYTEENABLE[22],f2h_sdram0_BYTEENABLE[21],f2h_sdram0_BYTEENABLE[20],f2h_sdram0_BYTEENABLE[19],f2h_sdram0_BYTEENABLE[18],f2h_sdram0_BYTEENABLE[17],f2h_sdram0_BYTEENABLE[16],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_sdram0_WRITEDATA[191],
f2h_sdram0_WRITEDATA[190],f2h_sdram0_WRITEDATA[189],f2h_sdram0_WRITEDATA[188],f2h_sdram0_WRITEDATA[187],f2h_sdram0_WRITEDATA[186],f2h_sdram0_WRITEDATA[185],f2h_sdram0_WRITEDATA[184],f2h_sdram0_WRITEDATA[183],f2h_sdram0_WRITEDATA[182],f2h_sdram0_WRITEDATA[181],f2h_sdram0_WRITEDATA[180],f2h_sdram0_WRITEDATA[179],
f2h_sdram0_WRITEDATA[178],f2h_sdram0_WRITEDATA[177],f2h_sdram0_WRITEDATA[176],f2h_sdram0_WRITEDATA[175],f2h_sdram0_WRITEDATA[174],f2h_sdram0_WRITEDATA[173],f2h_sdram0_WRITEDATA[172],f2h_sdram0_WRITEDATA[171],f2h_sdram0_WRITEDATA[170],f2h_sdram0_WRITEDATA[169],f2h_sdram0_WRITEDATA[168],f2h_sdram0_WRITEDATA[167],
f2h_sdram0_WRITEDATA[166],f2h_sdram0_WRITEDATA[165],f2h_sdram0_WRITEDATA[164],f2h_sdram0_WRITEDATA[163],f2h_sdram0_WRITEDATA[162],f2h_sdram0_WRITEDATA[161],f2h_sdram0_WRITEDATA[160],f2h_sdram0_WRITEDATA[159],f2h_sdram0_WRITEDATA[158],f2h_sdram0_WRITEDATA[157],f2h_sdram0_WRITEDATA[156],f2h_sdram0_WRITEDATA[155],
f2h_sdram0_WRITEDATA[154],f2h_sdram0_WRITEDATA[153],f2h_sdram0_WRITEDATA[152],f2h_sdram0_WRITEDATA[151],f2h_sdram0_WRITEDATA[150],f2h_sdram0_WRITEDATA[149],f2h_sdram0_WRITEDATA[148],f2h_sdram0_WRITEDATA[147],f2h_sdram0_WRITEDATA[146],f2h_sdram0_WRITEDATA[145],f2h_sdram0_WRITEDATA[144],f2h_sdram0_WRITEDATA[143],
f2h_sdram0_WRITEDATA[142],f2h_sdram0_WRITEDATA[141],f2h_sdram0_WRITEDATA[140],f2h_sdram0_WRITEDATA[139],f2h_sdram0_WRITEDATA[138],f2h_sdram0_WRITEDATA[137],f2h_sdram0_WRITEDATA[136],f2h_sdram0_WRITEDATA[135],f2h_sdram0_WRITEDATA[134],f2h_sdram0_WRITEDATA[133],f2h_sdram0_WRITEDATA[132],f2h_sdram0_WRITEDATA[131],
f2h_sdram0_WRITEDATA[130],f2h_sdram0_WRITEDATA[129],f2h_sdram0_WRITEDATA[128]}),
	.wr_data_3({gnd,gnd,f2h_sdram0_BYTEENABLE[31],f2h_sdram0_BYTEENABLE[30],f2h_sdram0_BYTEENABLE[29],f2h_sdram0_BYTEENABLE[28],f2h_sdram0_BYTEENABLE[27],f2h_sdram0_BYTEENABLE[26],f2h_sdram0_BYTEENABLE[25],f2h_sdram0_BYTEENABLE[24],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,f2h_sdram0_WRITEDATA[255],
f2h_sdram0_WRITEDATA[254],f2h_sdram0_WRITEDATA[253],f2h_sdram0_WRITEDATA[252],f2h_sdram0_WRITEDATA[251],f2h_sdram0_WRITEDATA[250],f2h_sdram0_WRITEDATA[249],f2h_sdram0_WRITEDATA[248],f2h_sdram0_WRITEDATA[247],f2h_sdram0_WRITEDATA[246],f2h_sdram0_WRITEDATA[245],f2h_sdram0_WRITEDATA[244],f2h_sdram0_WRITEDATA[243],
f2h_sdram0_WRITEDATA[242],f2h_sdram0_WRITEDATA[241],f2h_sdram0_WRITEDATA[240],f2h_sdram0_WRITEDATA[239],f2h_sdram0_WRITEDATA[238],f2h_sdram0_WRITEDATA[237],f2h_sdram0_WRITEDATA[236],f2h_sdram0_WRITEDATA[235],f2h_sdram0_WRITEDATA[234],f2h_sdram0_WRITEDATA[233],f2h_sdram0_WRITEDATA[232],f2h_sdram0_WRITEDATA[231],
f2h_sdram0_WRITEDATA[230],f2h_sdram0_WRITEDATA[229],f2h_sdram0_WRITEDATA[228],f2h_sdram0_WRITEDATA[227],f2h_sdram0_WRITEDATA[226],f2h_sdram0_WRITEDATA[225],f2h_sdram0_WRITEDATA[224],f2h_sdram0_WRITEDATA[223],f2h_sdram0_WRITEDATA[222],f2h_sdram0_WRITEDATA[221],f2h_sdram0_WRITEDATA[220],f2h_sdram0_WRITEDATA[219],
f2h_sdram0_WRITEDATA[218],f2h_sdram0_WRITEDATA[217],f2h_sdram0_WRITEDATA[216],f2h_sdram0_WRITEDATA[215],f2h_sdram0_WRITEDATA[214],f2h_sdram0_WRITEDATA[213],f2h_sdram0_WRITEDATA[212],f2h_sdram0_WRITEDATA[211],f2h_sdram0_WRITEDATA[210],f2h_sdram0_WRITEDATA[209],f2h_sdram0_WRITEDATA[208],f2h_sdram0_WRITEDATA[207],
f2h_sdram0_WRITEDATA[206],f2h_sdram0_WRITEDATA[205],f2h_sdram0_WRITEDATA[204],f2h_sdram0_WRITEDATA[203],f2h_sdram0_WRITEDATA[202],f2h_sdram0_WRITEDATA[201],f2h_sdram0_WRITEDATA[200],f2h_sdram0_WRITEDATA[199],f2h_sdram0_WRITEDATA[198],f2h_sdram0_WRITEDATA[197],f2h_sdram0_WRITEDATA[196],f2h_sdram0_WRITEDATA[195],
f2h_sdram0_WRITEDATA[194],f2h_sdram0_WRITEDATA[193],f2h_sdram0_WRITEDATA[192]}),
	.cmd_ready_0(f2h_sdram0_WAITREQUEST[0]),
	.cmd_ready_1(),
	.cmd_ready_2(),
	.cmd_ready_3(),
	.cmd_ready_4(),
	.cmd_ready_5(),
	.rd_valid_0(),
	.rd_valid_1(),
	.rd_valid_2(),
	.rd_valid_3(f2h_sdram0_READDATAVALID[0]),
	.wr_ready_0(),
	.wr_ready_1(),
	.wr_ready_2(),
	.wr_ready_3(),
	.wrack_valid_0(),
	.wrack_valid_1(),
	.wrack_valid_2(),
	.wrack_valid_3(),
	.wrack_valid_4(),
	.wrack_valid_5(),
	.bonding_out_1(f2sdram_BONDING_OUT_1_bus),
	.bonding_out_2(),
	.rd_data_0(f2sdram_RD_DATA_0_bus),
	.rd_data_1(f2sdram_RD_DATA_1_bus),
	.rd_data_2(f2sdram_RD_DATA_2_bus),
	.rd_data_3(f2sdram_RD_DATA_3_bus),
	.wrack_data_0(),
	.wrack_data_1(),
	.wrack_data_2(),
	.wrack_data_3(),
	.wrack_data_4(),
	.wrack_data_5());

cyclonev_lcell_comb \intermediate[12] (
	.dataa(!f2h_sdram0_READ[0]),
	.datab(!f2h_sdram0_WRITE[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\intermediate[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \intermediate[12] .extended_lut = "off";
defparam \intermediate[12] .lut_mask = 64'h7777777777777777;
defparam \intermediate[12] .shared_arith = "off";

cyclonev_hps_interface_dbg_apb debug_apb(
	.p_slv_err(gnd),
	.p_ready(gnd),
	.p_clk(gnd),
	.p_clk_en(gnd),
	.dbg_apb_disable(gnd),
	.p_rdata(32'b00000000000000000000000000000000),
	.p_addr_31(\debug_apb~O_P_ADDR_31 ),
	.p_write(),
	.p_sel(),
	.p_enable(),
	.p_reset_n(),
	.p_addr(),
	.p_wdata());
defparam debug_apb.dummy_param = 256;

cyclonev_hps_interface_stm_event stm_event(
	.stm_event({f2h_stm_hwevents[27],f2h_stm_hwevents[26],f2h_stm_hwevents[25],f2h_stm_hwevents[24],f2h_stm_hwevents[23],f2h_stm_hwevents[22],f2h_stm_hwevents[21],f2h_stm_hwevents[20],f2h_stm_hwevents[19],f2h_stm_hwevents[18],f2h_stm_hwevents[17],f2h_stm_hwevents[16],f2h_stm_hwevents[15],f2h_stm_hwevents[14],f2h_stm_hwevents[13],f2h_stm_hwevents[12],
f2h_stm_hwevents[11],f2h_stm_hwevents[10],f2h_stm_hwevents[9],f2h_stm_hwevents[8],f2h_stm_hwevents[7],f2h_stm_hwevents[6],f2h_stm_hwevents[5],f2h_stm_hwevents[4],f2h_stm_hwevents[3],f2h_stm_hwevents[2],f2h_stm_hwevents[1],f2h_stm_hwevents[0]}),
	.fake_dout(\stm_event~fake_dout ));

cyclonev_hps_interface_tpiu_trace tpiu(
	.traceclk_ctl(vcc),
	.traceclkin(gnd),
	.traceclk(),
	.trace_data(tpiu_TRACE_DATA_bus));

cyclonev_hps_interface_boot_from_fpga boot_from_fpga(
	.boot_from_fpga_on_failure(gnd),
	.boot_from_fpga_ready(gnd),
	.bsel_en(gnd),
	.csel_en(gnd),
	.bsel({gnd,gnd,vcc}),
	.csel({gnd,vcc}),
	.fake_dout(\boot_from_fpga~fake_dout ));

cyclonev_hps_interface_fpga2hps fpga2hps(
	.arvalid(gnd),
	.awvalid(gnd),
	.bready(gnd),
	.clk(h2f_lw_axi_clk[0]),
	.rready(gnd),
	.wlast(gnd),
	.wvalid(gnd),
	.araddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arburst({gnd,gnd}),
	.arcache({gnd,gnd,gnd,gnd}),
	.arid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arlen({gnd,gnd,gnd,gnd}),
	.arlock({gnd,gnd}),
	.arprot({gnd,gnd,gnd}),
	.arsize({gnd,gnd,gnd}),
	.aruser({gnd,gnd,gnd,gnd,gnd}),
	.awaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awburst({gnd,gnd}),
	.awcache({gnd,gnd,gnd,gnd}),
	.awid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.awlen({gnd,gnd,gnd,gnd}),
	.awlock({gnd,gnd}),
	.awprot({gnd,gnd,gnd}),
	.awsize({gnd,gnd,gnd}),
	.awuser({gnd,gnd,gnd,gnd,gnd}),
	.port_size_config({gnd,gnd}),
	.wdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.wstrb({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.arready(\f2h_ARREADY[0] ),
	.awready(),
	.bvalid(),
	.rlast(),
	.rvalid(),
	.wready(),
	.bid(),
	.bresp(),
	.rdata(),
	.rid(),
	.rresp());
defparam fpga2hps.data_width = 32;

cyclonev_hps_interface_hps2fpga hps2fpga(
	.arready(gnd),
	.awready(gnd),
	.bvalid(gnd),
	.clk(h2f_lw_axi_clk[0]),
	.rlast(gnd),
	.rvalid(gnd),
	.wready(gnd),
	.bid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.bresp({gnd,gnd}),
	.port_size_config({gnd,gnd}),
	.rdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rid({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.rresp({gnd,gnd}),
	.arvalid(),
	.awvalid(),
	.bready(),
	.rready(),
	.wlast(),
	.wvalid(),
	.araddr(hps2fpga_ARADDR_bus),
	.arburst(),
	.arcache(),
	.arid(),
	.arlen(),
	.arlock(),
	.arprot(),
	.arsize(),
	.awaddr(),
	.awburst(),
	.awcache(),
	.awid(),
	.awlen(),
	.awlock(),
	.awprot(),
	.awsize(),
	.wdata(),
	.wid(),
	.wstrb());
defparam hps2fpga.data_width = 32;

endmodule

module terminal_qsys_terminal_qsys_hps_hps_io (
	emac1_inst,
	emac1_inst1,
	intermediate_0,
	intermediate_1,
	emac1_inst2,
	emac1_inst3,
	emac1_inst4,
	emac1_inst5,
	emac1_inst6,
	sdio_inst,
	intermediate_2,
	intermediate_3,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_10,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	intermediate_11,
	uart0_inst,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_hps_io_hps_io_emac1_inst_RXD0,
	hps_hps_io_hps_io_emac1_inst_RXD1,
	hps_hps_io_hps_io_emac1_inst_RXD2,
	hps_hps_io_hps_io_emac1_inst_RXD3,
	hps_hps_io_hps_io_emac1_inst_RX_CLK,
	hps_hps_io_hps_io_emac1_inst_RX_CTL,
	hps_hps_io_hps_io_uart0_inst_RX,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	emac1_inst;
output 	emac1_inst1;
output 	intermediate_0;
output 	intermediate_1;
output 	emac1_inst2;
output 	emac1_inst3;
output 	emac1_inst4;
output 	emac1_inst5;
output 	emac1_inst6;
output 	sdio_inst;
output 	intermediate_2;
output 	intermediate_3;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_10;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	intermediate_11;
output 	uart0_inst;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	hps_hps_io_hps_io_emac1_inst_RXD0;
input 	hps_hps_io_hps_io_emac1_inst_RXD1;
input 	hps_hps_io_hps_io_emac1_inst_RXD2;
input 	hps_hps_io_hps_io_emac1_inst_RXD3;
input 	hps_hps_io_hps_io_emac1_inst_RX_CLK;
input 	hps_hps_io_hps_io_emac1_inst_RX_CTL;
input 	hps_hps_io_hps_io_uart0_inst_RX;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_terminal_qsys_hps_hps_io_border border(
	.hps_io_emac1_inst_TX_CLK({emac1_inst}),
	.hps_io_emac1_inst_TX_CTL({emac1_inst1}),
	.intermediate_0(intermediate_0),
	.intermediate_1(intermediate_1),
	.hps_io_emac1_inst_MDC({emac1_inst2}),
	.hps_io_emac1_inst_TXD0({emac1_inst3}),
	.hps_io_emac1_inst_TXD1({emac1_inst4}),
	.hps_io_emac1_inst_TXD2({emac1_inst5}),
	.hps_io_emac1_inst_TXD3({emac1_inst6}),
	.hps_io_sdio_inst_CLK({sdio_inst}),
	.intermediate_2(intermediate_2),
	.intermediate_3(intermediate_3),
	.intermediate_4(intermediate_4),
	.intermediate_6(intermediate_6),
	.intermediate_8(intermediate_8),
	.intermediate_10(intermediate_10),
	.intermediate_5(intermediate_5),
	.intermediate_7(intermediate_7),
	.intermediate_9(intermediate_9),
	.intermediate_11(intermediate_11),
	.hps_io_uart0_inst_TX({uart0_inst}),
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.hps_io_emac1_inst_MDIO_0(hps_io_emac1_inst_MDIO_0),
	.hps_io_sdio_inst_CMD_0(hps_io_sdio_inst_CMD_0),
	.hps_io_sdio_inst_D0_0(hps_io_sdio_inst_D0_0),
	.hps_io_sdio_inst_D1_0(hps_io_sdio_inst_D1_0),
	.hps_io_sdio_inst_D2_0(hps_io_sdio_inst_D2_0),
	.hps_io_sdio_inst_D3_0(hps_io_sdio_inst_D3_0),
	.hps_io_emac1_inst_RXD0({hps_hps_io_hps_io_emac1_inst_RXD0}),
	.hps_io_emac1_inst_RXD1({hps_hps_io_hps_io_emac1_inst_RXD1}),
	.hps_io_emac1_inst_RXD2({hps_hps_io_hps_io_emac1_inst_RXD2}),
	.hps_io_emac1_inst_RXD3({hps_hps_io_hps_io_emac1_inst_RXD3}),
	.hps_io_emac1_inst_RX_CLK({hps_hps_io_hps_io_emac1_inst_RX_CLK}),
	.hps_io_emac1_inst_RX_CTL({hps_hps_io_hps_io_emac1_inst_RX_CTL}),
	.hps_io_uart0_inst_RX({hps_hps_io_hps_io_uart0_inst_RX}),
	.memory_oct_rzqin(memory_oct_rzqin));

endmodule

module terminal_qsys_terminal_qsys_hps_hps_io_border (
	hps_io_emac1_inst_TX_CLK,
	hps_io_emac1_inst_TX_CTL,
	intermediate_0,
	intermediate_1,
	hps_io_emac1_inst_MDC,
	hps_io_emac1_inst_TXD0,
	hps_io_emac1_inst_TXD1,
	hps_io_emac1_inst_TXD2,
	hps_io_emac1_inst_TXD3,
	hps_io_sdio_inst_CLK,
	intermediate_2,
	intermediate_3,
	intermediate_4,
	intermediate_6,
	intermediate_8,
	intermediate_10,
	intermediate_5,
	intermediate_7,
	intermediate_9,
	intermediate_11,
	hps_io_uart0_inst_TX,
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	hps_io_emac1_inst_MDIO_0,
	hps_io_sdio_inst_CMD_0,
	hps_io_sdio_inst_D0_0,
	hps_io_sdio_inst_D1_0,
	hps_io_sdio_inst_D2_0,
	hps_io_sdio_inst_D3_0,
	hps_io_emac1_inst_RXD0,
	hps_io_emac1_inst_RXD1,
	hps_io_emac1_inst_RXD2,
	hps_io_emac1_inst_RXD3,
	hps_io_emac1_inst_RX_CLK,
	hps_io_emac1_inst_RX_CTL,
	hps_io_uart0_inst_RX,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[0:0] hps_io_emac1_inst_TX_CLK;
output 	[0:0] hps_io_emac1_inst_TX_CTL;
output 	intermediate_0;
output 	intermediate_1;
output 	[0:0] hps_io_emac1_inst_MDC;
output 	[0:0] hps_io_emac1_inst_TXD0;
output 	[0:0] hps_io_emac1_inst_TXD1;
output 	[0:0] hps_io_emac1_inst_TXD2;
output 	[0:0] hps_io_emac1_inst_TXD3;
output 	[0:0] hps_io_sdio_inst_CLK;
output 	intermediate_2;
output 	intermediate_3;
output 	intermediate_4;
output 	intermediate_6;
output 	intermediate_8;
output 	intermediate_10;
output 	intermediate_5;
output 	intermediate_7;
output 	intermediate_9;
output 	intermediate_11;
output 	[0:0] hps_io_uart0_inst_TX;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	hps_io_emac1_inst_MDIO_0;
input 	hps_io_sdio_inst_CMD_0;
input 	hps_io_sdio_inst_D0_0;
input 	hps_io_sdio_inst_D1_0;
input 	hps_io_sdio_inst_D2_0;
input 	hps_io_sdio_inst_D3_0;
input 	[0:0] hps_io_emac1_inst_RXD0;
input 	[0:0] hps_io_emac1_inst_RXD1;
input 	[0:0] hps_io_emac1_inst_RXD2;
input 	[0:0] hps_io_emac1_inst_RXD3;
input 	[0:0] hps_io_emac1_inst_RX_CLK;
input 	[0:0] hps_io_emac1_inst_RX_CTL;
input 	[0:0] hps_io_uart0_inst_RX;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sdio_inst~O_SDMMC_PWR_EN ;
wire \uart0_inst~UARTRTSN ;
wire \~GND~combout ;

wire [3:0] emac1_inst_EMAC_PHY_TXD_bus;
wire [7:0] sdio_inst_SDMMC_DATA_OE_bus;
wire [7:0] sdio_inst_SDMMC_DATA_O_bus;

assign hps_io_emac1_inst_TXD0[0] = emac1_inst_EMAC_PHY_TXD_bus[0];
assign hps_io_emac1_inst_TXD1[0] = emac1_inst_EMAC_PHY_TXD_bus[1];
assign hps_io_emac1_inst_TXD2[0] = emac1_inst_EMAC_PHY_TXD_bus[2];
assign hps_io_emac1_inst_TXD3[0] = emac1_inst_EMAC_PHY_TXD_bus[3];

assign intermediate_5 = sdio_inst_SDMMC_DATA_OE_bus[0];
assign intermediate_7 = sdio_inst_SDMMC_DATA_OE_bus[1];
assign intermediate_9 = sdio_inst_SDMMC_DATA_OE_bus[2];
assign intermediate_11 = sdio_inst_SDMMC_DATA_OE_bus[3];

assign intermediate_4 = sdio_inst_SDMMC_DATA_O_bus[0];
assign intermediate_6 = sdio_inst_SDMMC_DATA_O_bus[1];
assign intermediate_8 = sdio_inst_SDMMC_DATA_O_bus[2];
assign intermediate_10 = sdio_inst_SDMMC_DATA_O_bus[3];

terminal_qsys_hps_sdram hps_sdram_inst(
	.parallelterminationcontrol_0(parallelterminationcontrol_0),
	.parallelterminationcontrol_1(parallelterminationcontrol_1),
	.parallelterminationcontrol_2(parallelterminationcontrol_2),
	.parallelterminationcontrol_3(parallelterminationcontrol_3),
	.parallelterminationcontrol_4(parallelterminationcontrol_4),
	.parallelterminationcontrol_5(parallelterminationcontrol_5),
	.parallelterminationcontrol_6(parallelterminationcontrol_6),
	.parallelterminationcontrol_7(parallelterminationcontrol_7),
	.parallelterminationcontrol_8(parallelterminationcontrol_8),
	.parallelterminationcontrol_9(parallelterminationcontrol_9),
	.parallelterminationcontrol_10(parallelterminationcontrol_10),
	.parallelterminationcontrol_11(parallelterminationcontrol_11),
	.parallelterminationcontrol_12(parallelterminationcontrol_12),
	.parallelterminationcontrol_13(parallelterminationcontrol_13),
	.parallelterminationcontrol_14(parallelterminationcontrol_14),
	.parallelterminationcontrol_15(parallelterminationcontrol_15),
	.seriesterminationcontrol_0(seriesterminationcontrol_0),
	.seriesterminationcontrol_1(seriesterminationcontrol_1),
	.seriesterminationcontrol_2(seriesterminationcontrol_2),
	.seriesterminationcontrol_3(seriesterminationcontrol_3),
	.seriesterminationcontrol_4(seriesterminationcontrol_4),
	.seriesterminationcontrol_5(seriesterminationcontrol_5),
	.seriesterminationcontrol_6(seriesterminationcontrol_6),
	.seriesterminationcontrol_7(seriesterminationcontrol_7),
	.seriesterminationcontrol_8(seriesterminationcontrol_8),
	.seriesterminationcontrol_9(seriesterminationcontrol_9),
	.seriesterminationcontrol_10(seriesterminationcontrol_10),
	.seriesterminationcontrol_11(seriesterminationcontrol_11),
	.seriesterminationcontrol_12(seriesterminationcontrol_12),
	.seriesterminationcontrol_13(seriesterminationcontrol_13),
	.seriesterminationcontrol_14(seriesterminationcontrol_14),
	.seriesterminationcontrol_15(seriesterminationcontrol_15),
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.GND_port(\~GND~combout ),
	.memory_oct_rzqin(memory_oct_rzqin));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_hps_peripheral_emac emac1_inst(
	.emac_clk_rx(hps_io_emac1_inst_RX_CLK[0]),
	.emac_phy_rxdv(hps_io_emac1_inst_RX_CTL[0]),
	.emac_gmii_mdo_i(hps_io_emac1_inst_MDIO_0),
	.emac_phy_rxd({hps_io_emac1_inst_RXD3[0],hps_io_emac1_inst_RXD2[0],hps_io_emac1_inst_RXD1[0],hps_io_emac1_inst_RXD0[0]}),
	.emac_clk_tx(hps_io_emac1_inst_TX_CLK[0]),
	.emac_phy_tx_oe(hps_io_emac1_inst_TX_CTL[0]),
	.emac_gmii_mdo_o(intermediate_0),
	.emac_gmii_mdo_oe(intermediate_1),
	.emac_gmii_mdc(hps_io_emac1_inst_MDC[0]),
	.emac_phy_txd(emac1_inst_EMAC_PHY_TXD_bus));
defparam emac1_inst.dummy_param = 256;

cyclonev_hps_peripheral_sdmmc sdio_inst(
	.sdmmc_fb_clk(gnd),
	.sdmmc_cmd_i(hps_io_sdio_inst_CMD_0),
	.sdmmc_data_i({gnd,gnd,gnd,gnd,hps_io_sdio_inst_D3_0,hps_io_sdio_inst_D2_0,hps_io_sdio_inst_D1_0,hps_io_sdio_inst_D0_0}),
	.sdmmc_pwr_en(\sdio_inst~O_SDMMC_PWR_EN ),
	.sdmmc_cclk(hps_io_sdio_inst_CLK[0]),
	.sdmmc_cmd_o(intermediate_2),
	.sdmmc_cmd_oe(intermediate_3),
	.sdmmc_data_o(sdio_inst_SDMMC_DATA_O_bus),
	.sdmmc_data_oe(sdio_inst_SDMMC_DATA_OE_bus));
defparam sdio_inst.dummy_param = 256;

cyclonev_hps_peripheral_uart uart0_inst(
	.uart_cts_n(gnd),
	.uart_rxd(hps_io_uart0_inst_RX[0]),
	.uart_rts_n(\uart0_inst~UARTRTSN ),
	.uart_txd(hps_io_uart0_inst_TX[0]));
defparam uart0_inst.dummy_param = 256;

endmodule

module terminal_qsys_hps_sdram (
	parallelterminationcontrol_0,
	parallelterminationcontrol_1,
	parallelterminationcontrol_2,
	parallelterminationcontrol_3,
	parallelterminationcontrol_4,
	parallelterminationcontrol_5,
	parallelterminationcontrol_6,
	parallelterminationcontrol_7,
	parallelterminationcontrol_8,
	parallelterminationcontrol_9,
	parallelterminationcontrol_10,
	parallelterminationcontrol_11,
	parallelterminationcontrol_12,
	parallelterminationcontrol_13,
	parallelterminationcontrol_14,
	parallelterminationcontrol_15,
	seriesterminationcontrol_0,
	seriesterminationcontrol_1,
	seriesterminationcontrol_2,
	seriesterminationcontrol_3,
	seriesterminationcontrol_4,
	seriesterminationcontrol_5,
	seriesterminationcontrol_6,
	seriesterminationcontrol_7,
	seriesterminationcontrol_8,
	seriesterminationcontrol_9,
	seriesterminationcontrol_10,
	seriesterminationcontrol_11,
	seriesterminationcontrol_12,
	seriesterminationcontrol_13,
	seriesterminationcontrol_14,
	seriesterminationcontrol_15,
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	GND_port,
	memory_oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	parallelterminationcontrol_0;
output 	parallelterminationcontrol_1;
output 	parallelterminationcontrol_2;
output 	parallelterminationcontrol_3;
output 	parallelterminationcontrol_4;
output 	parallelterminationcontrol_5;
output 	parallelterminationcontrol_6;
output 	parallelterminationcontrol_7;
output 	parallelterminationcontrol_8;
output 	parallelterminationcontrol_9;
output 	parallelterminationcontrol_10;
output 	parallelterminationcontrol_11;
output 	parallelterminationcontrol_12;
output 	parallelterminationcontrol_13;
output 	parallelterminationcontrol_14;
output 	parallelterminationcontrol_15;
output 	seriesterminationcontrol_0;
output 	seriesterminationcontrol_1;
output 	seriesterminationcontrol_2;
output 	seriesterminationcontrol_3;
output 	seriesterminationcontrol_4;
output 	seriesterminationcontrol_5;
output 	seriesterminationcontrol_6;
output 	seriesterminationcontrol_7;
output 	seriesterminationcontrol_8;
output 	seriesterminationcontrol_9;
output 	seriesterminationcontrol_10;
output 	seriesterminationcontrol_11;
output 	seriesterminationcontrol_12;
output 	seriesterminationcontrol_13;
output 	seriesterminationcontrol_14;
output 	seriesterminationcontrol_15;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	GND_port;
input 	memory_oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pll|afi_clk ;
wire \pll|pll_write_clk ;
wire \p0|umemphy|afi_cal_fail ;
wire \p0|umemphy|afi_cal_success ;
wire \p0|umemphy|afi_rdata_valid[0] ;
wire \p0|umemphy|ctl_reset_n ;
wire \p0|umemphy|afi_rdata[0] ;
wire \p0|umemphy|afi_rdata[1] ;
wire \p0|umemphy|afi_rdata[2] ;
wire \p0|umemphy|afi_rdata[3] ;
wire \p0|umemphy|afi_rdata[4] ;
wire \p0|umemphy|afi_rdata[5] ;
wire \p0|umemphy|afi_rdata[6] ;
wire \p0|umemphy|afi_rdata[7] ;
wire \p0|umemphy|afi_rdata[8] ;
wire \p0|umemphy|afi_rdata[9] ;
wire \p0|umemphy|afi_rdata[10] ;
wire \p0|umemphy|afi_rdata[11] ;
wire \p0|umemphy|afi_rdata[12] ;
wire \p0|umemphy|afi_rdata[13] ;
wire \p0|umemphy|afi_rdata[14] ;
wire \p0|umemphy|afi_rdata[15] ;
wire \p0|umemphy|afi_rdata[16] ;
wire \p0|umemphy|afi_rdata[17] ;
wire \p0|umemphy|afi_rdata[18] ;
wire \p0|umemphy|afi_rdata[19] ;
wire \p0|umemphy|afi_rdata[20] ;
wire \p0|umemphy|afi_rdata[21] ;
wire \p0|umemphy|afi_rdata[22] ;
wire \p0|umemphy|afi_rdata[23] ;
wire \p0|umemphy|afi_rdata[24] ;
wire \p0|umemphy|afi_rdata[25] ;
wire \p0|umemphy|afi_rdata[26] ;
wire \p0|umemphy|afi_rdata[27] ;
wire \p0|umemphy|afi_rdata[28] ;
wire \p0|umemphy|afi_rdata[29] ;
wire \p0|umemphy|afi_rdata[30] ;
wire \p0|umemphy|afi_rdata[31] ;
wire \p0|umemphy|afi_rdata[32] ;
wire \p0|umemphy|afi_rdata[33] ;
wire \p0|umemphy|afi_rdata[34] ;
wire \p0|umemphy|afi_rdata[35] ;
wire \p0|umemphy|afi_rdata[36] ;
wire \p0|umemphy|afi_rdata[37] ;
wire \p0|umemphy|afi_rdata[38] ;
wire \p0|umemphy|afi_rdata[39] ;
wire \p0|umemphy|afi_rdata[40] ;
wire \p0|umemphy|afi_rdata[41] ;
wire \p0|umemphy|afi_rdata[42] ;
wire \p0|umemphy|afi_rdata[43] ;
wire \p0|umemphy|afi_rdata[44] ;
wire \p0|umemphy|afi_rdata[45] ;
wire \p0|umemphy|afi_rdata[46] ;
wire \p0|umemphy|afi_rdata[47] ;
wire \p0|umemphy|afi_rdata[48] ;
wire \p0|umemphy|afi_rdata[49] ;
wire \p0|umemphy|afi_rdata[50] ;
wire \p0|umemphy|afi_rdata[51] ;
wire \p0|umemphy|afi_rdata[52] ;
wire \p0|umemphy|afi_rdata[53] ;
wire \p0|umemphy|afi_rdata[54] ;
wire \p0|umemphy|afi_rdata[55] ;
wire \p0|umemphy|afi_rdata[56] ;
wire \p0|umemphy|afi_rdata[57] ;
wire \p0|umemphy|afi_rdata[58] ;
wire \p0|umemphy|afi_rdata[59] ;
wire \p0|umemphy|afi_rdata[60] ;
wire \p0|umemphy|afi_rdata[61] ;
wire \p0|umemphy|afi_rdata[62] ;
wire \p0|umemphy|afi_rdata[63] ;
wire \p0|umemphy|afi_rdata[64] ;
wire \p0|umemphy|afi_rdata[65] ;
wire \p0|umemphy|afi_rdata[66] ;
wire \p0|umemphy|afi_rdata[67] ;
wire \p0|umemphy|afi_rdata[68] ;
wire \p0|umemphy|afi_rdata[69] ;
wire \p0|umemphy|afi_rdata[70] ;
wire \p0|umemphy|afi_rdata[71] ;
wire \p0|umemphy|afi_rdata[72] ;
wire \p0|umemphy|afi_rdata[73] ;
wire \p0|umemphy|afi_rdata[74] ;
wire \p0|umemphy|afi_rdata[75] ;
wire \p0|umemphy|afi_rdata[76] ;
wire \p0|umemphy|afi_rdata[77] ;
wire \p0|umemphy|afi_rdata[78] ;
wire \p0|umemphy|afi_rdata[79] ;
wire \p0|umemphy|afi_wlat[0] ;
wire \p0|umemphy|afi_wlat[1] ;
wire \p0|umemphy|afi_wlat[2] ;
wire \p0|umemphy|afi_wlat[3] ;
wire \c0|afi_cas_n[0] ;
wire \c0|afi_ras_n[0] ;
wire \c0|afi_rst_n[0] ;
wire \c0|afi_we_n[0] ;
wire \c0|afi_addr[0] ;
wire \c0|afi_addr[1] ;
wire \c0|afi_addr[2] ;
wire \c0|afi_addr[3] ;
wire \c0|afi_addr[4] ;
wire \c0|afi_addr[5] ;
wire \c0|afi_addr[6] ;
wire \c0|afi_addr[7] ;
wire \c0|afi_addr[8] ;
wire \c0|afi_addr[9] ;
wire \c0|afi_addr[10] ;
wire \c0|afi_addr[11] ;
wire \c0|afi_addr[12] ;
wire \c0|afi_addr[13] ;
wire \c0|afi_addr[14] ;
wire \c0|afi_addr[15] ;
wire \c0|afi_addr[16] ;
wire \c0|afi_addr[17] ;
wire \c0|afi_addr[18] ;
wire \c0|afi_addr[19] ;
wire \c0|afi_ba[0] ;
wire \c0|afi_ba[1] ;
wire \c0|afi_ba[2] ;
wire \c0|afi_cke[0] ;
wire \c0|afi_cke[1] ;
wire \c0|afi_cs_n[0] ;
wire \c0|afi_cs_n[1] ;
wire \c0|afi_dm_int[0] ;
wire \c0|afi_dm_int[1] ;
wire \c0|afi_dm_int[2] ;
wire \c0|afi_dm_int[3] ;
wire \c0|afi_dm_int[4] ;
wire \c0|afi_dm_int[5] ;
wire \c0|afi_dm_int[6] ;
wire \c0|afi_dm_int[7] ;
wire \c0|afi_dm_int[8] ;
wire \c0|afi_dm_int[9] ;
wire \c0|afi_dqs_burst[0] ;
wire \c0|afi_dqs_burst[1] ;
wire \c0|afi_dqs_burst[2] ;
wire \c0|afi_dqs_burst[3] ;
wire \c0|afi_dqs_burst[4] ;
wire \c0|afi_odt[0] ;
wire \c0|afi_odt[1] ;
wire \c0|afi_rdata_en[0] ;
wire \c0|afi_rdata_en[1] ;
wire \c0|afi_rdata_en[2] ;
wire \c0|afi_rdata_en[3] ;
wire \c0|afi_rdata_en[4] ;
wire \c0|afi_rdata_en_full[0] ;
wire \c0|afi_rdata_en_full[1] ;
wire \c0|afi_rdata_en_full[2] ;
wire \c0|afi_rdata_en_full[3] ;
wire \c0|afi_rdata_en_full[4] ;
wire \c0|afi_wdata_int[0] ;
wire \c0|afi_wdata_int[1] ;
wire \c0|afi_wdata_int[2] ;
wire \c0|afi_wdata_int[3] ;
wire \c0|afi_wdata_int[4] ;
wire \c0|afi_wdata_int[5] ;
wire \c0|afi_wdata_int[6] ;
wire \c0|afi_wdata_int[7] ;
wire \c0|afi_wdata_int[8] ;
wire \c0|afi_wdata_int[9] ;
wire \c0|afi_wdata_int[10] ;
wire \c0|afi_wdata_int[11] ;
wire \c0|afi_wdata_int[12] ;
wire \c0|afi_wdata_int[13] ;
wire \c0|afi_wdata_int[14] ;
wire \c0|afi_wdata_int[15] ;
wire \c0|afi_wdata_int[16] ;
wire \c0|afi_wdata_int[17] ;
wire \c0|afi_wdata_int[18] ;
wire \c0|afi_wdata_int[19] ;
wire \c0|afi_wdata_int[20] ;
wire \c0|afi_wdata_int[21] ;
wire \c0|afi_wdata_int[22] ;
wire \c0|afi_wdata_int[23] ;
wire \c0|afi_wdata_int[24] ;
wire \c0|afi_wdata_int[25] ;
wire \c0|afi_wdata_int[26] ;
wire \c0|afi_wdata_int[27] ;
wire \c0|afi_wdata_int[28] ;
wire \c0|afi_wdata_int[29] ;
wire \c0|afi_wdata_int[30] ;
wire \c0|afi_wdata_int[31] ;
wire \c0|afi_wdata_int[32] ;
wire \c0|afi_wdata_int[33] ;
wire \c0|afi_wdata_int[34] ;
wire \c0|afi_wdata_int[35] ;
wire \c0|afi_wdata_int[36] ;
wire \c0|afi_wdata_int[37] ;
wire \c0|afi_wdata_int[38] ;
wire \c0|afi_wdata_int[39] ;
wire \c0|afi_wdata_int[40] ;
wire \c0|afi_wdata_int[41] ;
wire \c0|afi_wdata_int[42] ;
wire \c0|afi_wdata_int[43] ;
wire \c0|afi_wdata_int[44] ;
wire \c0|afi_wdata_int[45] ;
wire \c0|afi_wdata_int[46] ;
wire \c0|afi_wdata_int[47] ;
wire \c0|afi_wdata_int[48] ;
wire \c0|afi_wdata_int[49] ;
wire \c0|afi_wdata_int[50] ;
wire \c0|afi_wdata_int[51] ;
wire \c0|afi_wdata_int[52] ;
wire \c0|afi_wdata_int[53] ;
wire \c0|afi_wdata_int[54] ;
wire \c0|afi_wdata_int[55] ;
wire \c0|afi_wdata_int[56] ;
wire \c0|afi_wdata_int[57] ;
wire \c0|afi_wdata_int[58] ;
wire \c0|afi_wdata_int[59] ;
wire \c0|afi_wdata_int[60] ;
wire \c0|afi_wdata_int[61] ;
wire \c0|afi_wdata_int[62] ;
wire \c0|afi_wdata_int[63] ;
wire \c0|afi_wdata_int[64] ;
wire \c0|afi_wdata_int[65] ;
wire \c0|afi_wdata_int[66] ;
wire \c0|afi_wdata_int[67] ;
wire \c0|afi_wdata_int[68] ;
wire \c0|afi_wdata_int[69] ;
wire \c0|afi_wdata_int[70] ;
wire \c0|afi_wdata_int[71] ;
wire \c0|afi_wdata_int[72] ;
wire \c0|afi_wdata_int[73] ;
wire \c0|afi_wdata_int[74] ;
wire \c0|afi_wdata_int[75] ;
wire \c0|afi_wdata_int[76] ;
wire \c0|afi_wdata_int[77] ;
wire \c0|afi_wdata_int[78] ;
wire \c0|afi_wdata_int[79] ;
wire \c0|afi_wdata_valid[0] ;
wire \c0|afi_wdata_valid[1] ;
wire \c0|afi_wdata_valid[2] ;
wire \c0|afi_wdata_valid[3] ;
wire \c0|afi_wdata_valid[4] ;
wire \c0|cfg_addlat_wire[0] ;
wire \c0|cfg_addlat_wire[1] ;
wire \c0|cfg_addlat_wire[2] ;
wire \c0|cfg_addlat_wire[3] ;
wire \c0|cfg_addlat_wire[4] ;
wire \c0|cfg_bankaddrwidth_wire[0] ;
wire \c0|cfg_bankaddrwidth_wire[1] ;
wire \c0|cfg_bankaddrwidth_wire[2] ;
wire \c0|cfg_caswrlat_wire[0] ;
wire \c0|cfg_caswrlat_wire[1] ;
wire \c0|cfg_caswrlat_wire[2] ;
wire \c0|cfg_caswrlat_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[0] ;
wire \c0|cfg_coladdrwidth_wire[1] ;
wire \c0|cfg_coladdrwidth_wire[2] ;
wire \c0|cfg_coladdrwidth_wire[3] ;
wire \c0|cfg_coladdrwidth_wire[4] ;
wire \c0|cfg_csaddrwidth_wire[0] ;
wire \c0|cfg_csaddrwidth_wire[1] ;
wire \c0|cfg_csaddrwidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[0] ;
wire \c0|cfg_devicewidth_wire[1] ;
wire \c0|cfg_devicewidth_wire[2] ;
wire \c0|cfg_devicewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[0] ;
wire \c0|cfg_interfacewidth_wire[1] ;
wire \c0|cfg_interfacewidth_wire[2] ;
wire \c0|cfg_interfacewidth_wire[3] ;
wire \c0|cfg_interfacewidth_wire[4] ;
wire \c0|cfg_interfacewidth_wire[5] ;
wire \c0|cfg_interfacewidth_wire[6] ;
wire \c0|cfg_interfacewidth_wire[7] ;
wire \c0|cfg_rowaddrwidth_wire[0] ;
wire \c0|cfg_rowaddrwidth_wire[1] ;
wire \c0|cfg_rowaddrwidth_wire[2] ;
wire \c0|cfg_rowaddrwidth_wire[3] ;
wire \c0|cfg_rowaddrwidth_wire[4] ;
wire \c0|cfg_tcl_wire[0] ;
wire \c0|cfg_tcl_wire[1] ;
wire \c0|cfg_tcl_wire[2] ;
wire \c0|cfg_tcl_wire[3] ;
wire \c0|cfg_tcl_wire[4] ;
wire \c0|cfg_tmrd_wire[0] ;
wire \c0|cfg_tmrd_wire[1] ;
wire \c0|cfg_tmrd_wire[2] ;
wire \c0|cfg_tmrd_wire[3] ;
wire \c0|cfg_trefi_wire[0] ;
wire \c0|cfg_trefi_wire[1] ;
wire \c0|cfg_trefi_wire[2] ;
wire \c0|cfg_trefi_wire[3] ;
wire \c0|cfg_trefi_wire[4] ;
wire \c0|cfg_trefi_wire[5] ;
wire \c0|cfg_trefi_wire[6] ;
wire \c0|cfg_trefi_wire[7] ;
wire \c0|cfg_trefi_wire[8] ;
wire \c0|cfg_trefi_wire[9] ;
wire \c0|cfg_trefi_wire[10] ;
wire \c0|cfg_trefi_wire[11] ;
wire \c0|cfg_trefi_wire[12] ;
wire \c0|cfg_trfc_wire[0] ;
wire \c0|cfg_trfc_wire[1] ;
wire \c0|cfg_trfc_wire[2] ;
wire \c0|cfg_trfc_wire[3] ;
wire \c0|cfg_trfc_wire[4] ;
wire \c0|cfg_trfc_wire[5] ;
wire \c0|cfg_trfc_wire[6] ;
wire \c0|cfg_trfc_wire[7] ;
wire \c0|cfg_twr_wire[0] ;
wire \c0|cfg_twr_wire[1] ;
wire \c0|cfg_twr_wire[2] ;
wire \c0|cfg_twr_wire[3] ;
wire \c0|afi_mem_clk_disable[0] ;
wire \c0|cfg_dramconfig_wire[0] ;
wire \c0|cfg_dramconfig_wire[1] ;
wire \c0|cfg_dramconfig_wire[2] ;
wire \c0|cfg_dramconfig_wire[3] ;
wire \c0|cfg_dramconfig_wire[4] ;
wire \c0|cfg_dramconfig_wire[5] ;
wire \c0|cfg_dramconfig_wire[6] ;
wire \c0|cfg_dramconfig_wire[7] ;
wire \c0|cfg_dramconfig_wire[8] ;
wire \c0|cfg_dramconfig_wire[9] ;
wire \c0|cfg_dramconfig_wire[10] ;
wire \c0|cfg_dramconfig_wire[11] ;
wire \c0|cfg_dramconfig_wire[12] ;
wire \c0|cfg_dramconfig_wire[13] ;
wire \c0|cfg_dramconfig_wire[14] ;
wire \c0|cfg_dramconfig_wire[15] ;
wire \c0|cfg_dramconfig_wire[16] ;
wire \c0|cfg_dramconfig_wire[17] ;
wire \c0|cfg_dramconfig_wire[18] ;
wire \c0|cfg_dramconfig_wire[19] ;
wire \c0|cfg_dramconfig_wire[20] ;
wire \p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ;
wire \dll|dll_delayctrl[0] ;
wire \dll|dll_delayctrl[1] ;
wire \dll|dll_delayctrl[2] ;
wire \dll|dll_delayctrl[3] ;
wire \dll|dll_delayctrl[4] ;
wire \dll|dll_delayctrl[5] ;
wire \dll|dll_delayctrl[6] ;


terminal_qsys_altera_mem_if_dll_cyclonev dll(
	.clk(\pll|pll_write_clk ),
	.dll_delayctrl({\dll|dll_delayctrl[6] ,\dll|dll_delayctrl[5] ,\dll|dll_delayctrl[4] ,\dll|dll_delayctrl[3] ,\dll|dll_delayctrl[2] ,\dll|dll_delayctrl[1] ,\dll|dll_delayctrl[0] }));

terminal_qsys_altera_mem_if_oct_cyclonev oct(
	.parallelterminationcontrol({parallelterminationcontrol_15,parallelterminationcontrol_14,parallelterminationcontrol_13,parallelterminationcontrol_12,parallelterminationcontrol_11,parallelterminationcontrol_10,parallelterminationcontrol_9,parallelterminationcontrol_8,
parallelterminationcontrol_7,parallelterminationcontrol_6,parallelterminationcontrol_5,parallelterminationcontrol_4,parallelterminationcontrol_3,parallelterminationcontrol_2,parallelterminationcontrol_1,parallelterminationcontrol_0}),
	.seriesterminationcontrol({seriesterminationcontrol_15,seriesterminationcontrol_14,seriesterminationcontrol_13,seriesterminationcontrol_12,seriesterminationcontrol_11,seriesterminationcontrol_10,seriesterminationcontrol_9,seriesterminationcontrol_8,seriesterminationcontrol_7,
seriesterminationcontrol_6,seriesterminationcontrol_5,seriesterminationcontrol_4,seriesterminationcontrol_3,seriesterminationcontrol_2,seriesterminationcontrol_1,seriesterminationcontrol_0}),
	.oct_rzqin(memory_oct_rzqin));

terminal_qsys_altera_mem_if_hard_memory_controller_top_cyclonev c0(
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid({\p0|umemphy|afi_rdata_valid[0] }),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata({\p0|umemphy|afi_rdata[79] ,\p0|umemphy|afi_rdata[78] ,\p0|umemphy|afi_rdata[77] ,\p0|umemphy|afi_rdata[76] ,\p0|umemphy|afi_rdata[75] ,\p0|umemphy|afi_rdata[74] ,\p0|umemphy|afi_rdata[73] ,\p0|umemphy|afi_rdata[72] ,\p0|umemphy|afi_rdata[71] ,
\p0|umemphy|afi_rdata[70] ,\p0|umemphy|afi_rdata[69] ,\p0|umemphy|afi_rdata[68] ,\p0|umemphy|afi_rdata[67] ,\p0|umemphy|afi_rdata[66] ,\p0|umemphy|afi_rdata[65] ,\p0|umemphy|afi_rdata[64] ,\p0|umemphy|afi_rdata[63] ,\p0|umemphy|afi_rdata[62] ,
\p0|umemphy|afi_rdata[61] ,\p0|umemphy|afi_rdata[60] ,\p0|umemphy|afi_rdata[59] ,\p0|umemphy|afi_rdata[58] ,\p0|umemphy|afi_rdata[57] ,\p0|umemphy|afi_rdata[56] ,\p0|umemphy|afi_rdata[55] ,\p0|umemphy|afi_rdata[54] ,\p0|umemphy|afi_rdata[53] ,
\p0|umemphy|afi_rdata[52] ,\p0|umemphy|afi_rdata[51] ,\p0|umemphy|afi_rdata[50] ,\p0|umemphy|afi_rdata[49] ,\p0|umemphy|afi_rdata[48] ,\p0|umemphy|afi_rdata[47] ,\p0|umemphy|afi_rdata[46] ,\p0|umemphy|afi_rdata[45] ,\p0|umemphy|afi_rdata[44] ,
\p0|umemphy|afi_rdata[43] ,\p0|umemphy|afi_rdata[42] ,\p0|umemphy|afi_rdata[41] ,\p0|umemphy|afi_rdata[40] ,\p0|umemphy|afi_rdata[39] ,\p0|umemphy|afi_rdata[38] ,\p0|umemphy|afi_rdata[37] ,\p0|umemphy|afi_rdata[36] ,\p0|umemphy|afi_rdata[35] ,
\p0|umemphy|afi_rdata[34] ,\p0|umemphy|afi_rdata[33] ,\p0|umemphy|afi_rdata[32] ,\p0|umemphy|afi_rdata[31] ,\p0|umemphy|afi_rdata[30] ,\p0|umemphy|afi_rdata[29] ,\p0|umemphy|afi_rdata[28] ,\p0|umemphy|afi_rdata[27] ,\p0|umemphy|afi_rdata[26] ,
\p0|umemphy|afi_rdata[25] ,\p0|umemphy|afi_rdata[24] ,\p0|umemphy|afi_rdata[23] ,\p0|umemphy|afi_rdata[22] ,\p0|umemphy|afi_rdata[21] ,\p0|umemphy|afi_rdata[20] ,\p0|umemphy|afi_rdata[19] ,\p0|umemphy|afi_rdata[18] ,\p0|umemphy|afi_rdata[17] ,
\p0|umemphy|afi_rdata[16] ,\p0|umemphy|afi_rdata[15] ,\p0|umemphy|afi_rdata[14] ,\p0|umemphy|afi_rdata[13] ,\p0|umemphy|afi_rdata[12] ,\p0|umemphy|afi_rdata[11] ,\p0|umemphy|afi_rdata[10] ,\p0|umemphy|afi_rdata[9] ,\p0|umemphy|afi_rdata[8] ,
\p0|umemphy|afi_rdata[7] ,\p0|umemphy|afi_rdata[6] ,\p0|umemphy|afi_rdata[5] ,\p0|umemphy|afi_rdata[4] ,\p0|umemphy|afi_rdata[3] ,\p0|umemphy|afi_rdata[2] ,\p0|umemphy|afi_rdata[1] ,\p0|umemphy|afi_rdata[0] }),
	.afi_wlat({\p0|umemphy|afi_wlat[3] ,\p0|umemphy|afi_wlat[2] ,\p0|umemphy|afi_wlat[1] ,\p0|umemphy|afi_wlat[0] }),
	.afi_cas_n({\c0|afi_cas_n[0] }),
	.afi_ras_n({\c0|afi_ras_n[0] }),
	.afi_rst_n({\c0|afi_rst_n[0] }),
	.afi_we_n({\c0|afi_we_n[0] }),
	.afi_addr({\c0|afi_addr[19] ,\c0|afi_addr[18] ,\c0|afi_addr[17] ,\c0|afi_addr[16] ,\c0|afi_addr[15] ,\c0|afi_addr[14] ,\c0|afi_addr[13] ,\c0|afi_addr[12] ,\c0|afi_addr[11] ,\c0|afi_addr[10] ,\c0|afi_addr[9] ,\c0|afi_addr[8] ,\c0|afi_addr[7] ,\c0|afi_addr[6] ,\c0|afi_addr[5] ,
\c0|afi_addr[4] ,\c0|afi_addr[3] ,\c0|afi_addr[2] ,\c0|afi_addr[1] ,\c0|afi_addr[0] }),
	.afi_ba({\c0|afi_ba[2] ,\c0|afi_ba[1] ,\c0|afi_ba[0] }),
	.afi_cke({\c0|afi_cke[1] ,\c0|afi_cke[0] }),
	.afi_cs_n({\c0|afi_cs_n[1] ,\c0|afi_cs_n[0] }),
	.afi_dm({\c0|afi_dm_int[9] ,\c0|afi_dm_int[8] ,\c0|afi_dm_int[7] ,\c0|afi_dm_int[6] ,\c0|afi_dm_int[5] ,\c0|afi_dm_int[4] ,\c0|afi_dm_int[3] ,\c0|afi_dm_int[2] ,\c0|afi_dm_int[1] ,\c0|afi_dm_int[0] }),
	.afi_dqs_burst({\c0|afi_dqs_burst[4] ,\c0|afi_dqs_burst[3] ,\c0|afi_dqs_burst[2] ,\c0|afi_dqs_burst[1] ,\c0|afi_dqs_burst[0] }),
	.afi_odt({\c0|afi_odt[1] ,\c0|afi_odt[0] }),
	.afi_rdata_en({\c0|afi_rdata_en[4] ,\c0|afi_rdata_en[3] ,\c0|afi_rdata_en[2] ,\c0|afi_rdata_en[1] ,\c0|afi_rdata_en[0] }),
	.afi_rdata_en_full({\c0|afi_rdata_en_full[4] ,\c0|afi_rdata_en_full[3] ,\c0|afi_rdata_en_full[2] ,\c0|afi_rdata_en_full[1] ,\c0|afi_rdata_en_full[0] }),
	.afi_wdata({\c0|afi_wdata_int[79] ,\c0|afi_wdata_int[78] ,\c0|afi_wdata_int[77] ,\c0|afi_wdata_int[76] ,\c0|afi_wdata_int[75] ,\c0|afi_wdata_int[74] ,\c0|afi_wdata_int[73] ,\c0|afi_wdata_int[72] ,\c0|afi_wdata_int[71] ,\c0|afi_wdata_int[70] ,\c0|afi_wdata_int[69] ,
\c0|afi_wdata_int[68] ,\c0|afi_wdata_int[67] ,\c0|afi_wdata_int[66] ,\c0|afi_wdata_int[65] ,\c0|afi_wdata_int[64] ,\c0|afi_wdata_int[63] ,\c0|afi_wdata_int[62] ,\c0|afi_wdata_int[61] ,\c0|afi_wdata_int[60] ,\c0|afi_wdata_int[59] ,\c0|afi_wdata_int[58] ,
\c0|afi_wdata_int[57] ,\c0|afi_wdata_int[56] ,\c0|afi_wdata_int[55] ,\c0|afi_wdata_int[54] ,\c0|afi_wdata_int[53] ,\c0|afi_wdata_int[52] ,\c0|afi_wdata_int[51] ,\c0|afi_wdata_int[50] ,\c0|afi_wdata_int[49] ,\c0|afi_wdata_int[48] ,\c0|afi_wdata_int[47] ,
\c0|afi_wdata_int[46] ,\c0|afi_wdata_int[45] ,\c0|afi_wdata_int[44] ,\c0|afi_wdata_int[43] ,\c0|afi_wdata_int[42] ,\c0|afi_wdata_int[41] ,\c0|afi_wdata_int[40] ,\c0|afi_wdata_int[39] ,\c0|afi_wdata_int[38] ,\c0|afi_wdata_int[37] ,\c0|afi_wdata_int[36] ,
\c0|afi_wdata_int[35] ,\c0|afi_wdata_int[34] ,\c0|afi_wdata_int[33] ,\c0|afi_wdata_int[32] ,\c0|afi_wdata_int[31] ,\c0|afi_wdata_int[30] ,\c0|afi_wdata_int[29] ,\c0|afi_wdata_int[28] ,\c0|afi_wdata_int[27] ,\c0|afi_wdata_int[26] ,\c0|afi_wdata_int[25] ,
\c0|afi_wdata_int[24] ,\c0|afi_wdata_int[23] ,\c0|afi_wdata_int[22] ,\c0|afi_wdata_int[21] ,\c0|afi_wdata_int[20] ,\c0|afi_wdata_int[19] ,\c0|afi_wdata_int[18] ,\c0|afi_wdata_int[17] ,\c0|afi_wdata_int[16] ,\c0|afi_wdata_int[15] ,\c0|afi_wdata_int[14] ,
\c0|afi_wdata_int[13] ,\c0|afi_wdata_int[12] ,\c0|afi_wdata_int[11] ,\c0|afi_wdata_int[10] ,\c0|afi_wdata_int[9] ,\c0|afi_wdata_int[8] ,\c0|afi_wdata_int[7] ,\c0|afi_wdata_int[6] ,\c0|afi_wdata_int[5] ,\c0|afi_wdata_int[4] ,\c0|afi_wdata_int[3] ,\c0|afi_wdata_int[2] ,
\c0|afi_wdata_int[1] ,\c0|afi_wdata_int[0] }),
	.afi_wdata_valid({\c0|afi_wdata_valid[4] ,\c0|afi_wdata_valid[3] ,\c0|afi_wdata_valid[2] ,\c0|afi_wdata_valid[1] ,\c0|afi_wdata_valid[0] }),
	.cfg_addlat({cfg_addlat_unconnected_wire_7,cfg_addlat_unconnected_wire_6,cfg_addlat_unconnected_wire_5,\c0|cfg_addlat_wire[4] ,\c0|cfg_addlat_wire[3] ,\c0|cfg_addlat_wire[2] ,\c0|cfg_addlat_wire[1] ,\c0|cfg_addlat_wire[0] }),
	.cfg_bankaddrwidth({cfg_bankaddrwidth_unconnected_wire_7,cfg_bankaddrwidth_unconnected_wire_6,cfg_bankaddrwidth_unconnected_wire_5,cfg_bankaddrwidth_unconnected_wire_4,cfg_bankaddrwidth_unconnected_wire_3,\c0|cfg_bankaddrwidth_wire[2] ,\c0|cfg_bankaddrwidth_wire[1] ,
\c0|cfg_bankaddrwidth_wire[0] }),
	.cfg_caswrlat({cfg_caswrlat_unconnected_wire_7,cfg_caswrlat_unconnected_wire_6,cfg_caswrlat_unconnected_wire_5,cfg_caswrlat_unconnected_wire_4,\c0|cfg_caswrlat_wire[3] ,\c0|cfg_caswrlat_wire[2] ,\c0|cfg_caswrlat_wire[1] ,\c0|cfg_caswrlat_wire[0] }),
	.cfg_coladdrwidth({cfg_coladdrwidth_unconnected_wire_7,cfg_coladdrwidth_unconnected_wire_6,cfg_coladdrwidth_unconnected_wire_5,\c0|cfg_coladdrwidth_wire[4] ,\c0|cfg_coladdrwidth_wire[3] ,\c0|cfg_coladdrwidth_wire[2] ,\c0|cfg_coladdrwidth_wire[1] ,\c0|cfg_coladdrwidth_wire[0] }),
	.cfg_csaddrwidth({cfg_csaddrwidth_unconnected_wire_7,cfg_csaddrwidth_unconnected_wire_6,cfg_csaddrwidth_unconnected_wire_5,cfg_csaddrwidth_unconnected_wire_4,cfg_csaddrwidth_unconnected_wire_3,\c0|cfg_csaddrwidth_wire[2] ,\c0|cfg_csaddrwidth_wire[1] ,\c0|cfg_csaddrwidth_wire[0] }),
	.cfg_devicewidth({cfg_devicewidth_unconnected_wire_7,cfg_devicewidth_unconnected_wire_6,cfg_devicewidth_unconnected_wire_5,cfg_devicewidth_unconnected_wire_4,\c0|cfg_devicewidth_wire[3] ,\c0|cfg_devicewidth_wire[2] ,\c0|cfg_devicewidth_wire[1] ,\c0|cfg_devicewidth_wire[0] }),
	.cfg_interfacewidth({\c0|cfg_interfacewidth_wire[7] ,\c0|cfg_interfacewidth_wire[6] ,\c0|cfg_interfacewidth_wire[5] ,\c0|cfg_interfacewidth_wire[4] ,\c0|cfg_interfacewidth_wire[3] ,\c0|cfg_interfacewidth_wire[2] ,\c0|cfg_interfacewidth_wire[1] ,\c0|cfg_interfacewidth_wire[0] }),
	.cfg_rowaddrwidth({cfg_rowaddrwidth_unconnected_wire_7,cfg_rowaddrwidth_unconnected_wire_6,cfg_rowaddrwidth_unconnected_wire_5,\c0|cfg_rowaddrwidth_wire[4] ,\c0|cfg_rowaddrwidth_wire[3] ,\c0|cfg_rowaddrwidth_wire[2] ,\c0|cfg_rowaddrwidth_wire[1] ,\c0|cfg_rowaddrwidth_wire[0] }),
	.cfg_tcl({cfg_tcl_unconnected_wire_7,cfg_tcl_unconnected_wire_6,cfg_tcl_unconnected_wire_5,\c0|cfg_tcl_wire[4] ,\c0|cfg_tcl_wire[3] ,\c0|cfg_tcl_wire[2] ,\c0|cfg_tcl_wire[1] ,\c0|cfg_tcl_wire[0] }),
	.cfg_tmrd({cfg_tmrd_unconnected_wire_7,cfg_tmrd_unconnected_wire_6,cfg_tmrd_unconnected_wire_5,cfg_tmrd_unconnected_wire_4,\c0|cfg_tmrd_wire[3] ,\c0|cfg_tmrd_wire[2] ,\c0|cfg_tmrd_wire[1] ,\c0|cfg_tmrd_wire[0] }),
	.cfg_trefi({cfg_trefi_unconnected_wire_15,cfg_trefi_unconnected_wire_14,cfg_trefi_unconnected_wire_13,\c0|cfg_trefi_wire[12] ,\c0|cfg_trefi_wire[11] ,\c0|cfg_trefi_wire[10] ,\c0|cfg_trefi_wire[9] ,\c0|cfg_trefi_wire[8] ,\c0|cfg_trefi_wire[7] ,\c0|cfg_trefi_wire[6] ,
\c0|cfg_trefi_wire[5] ,\c0|cfg_trefi_wire[4] ,\c0|cfg_trefi_wire[3] ,\c0|cfg_trefi_wire[2] ,\c0|cfg_trefi_wire[1] ,\c0|cfg_trefi_wire[0] }),
	.cfg_trfc({\c0|cfg_trfc_wire[7] ,\c0|cfg_trfc_wire[6] ,\c0|cfg_trfc_wire[5] ,\c0|cfg_trfc_wire[4] ,\c0|cfg_trfc_wire[3] ,\c0|cfg_trfc_wire[2] ,\c0|cfg_trfc_wire[1] ,\c0|cfg_trfc_wire[0] }),
	.cfg_twr({cfg_twr_unconnected_wire_7,cfg_twr_unconnected_wire_6,cfg_twr_unconnected_wire_5,cfg_twr_unconnected_wire_4,\c0|cfg_twr_wire[3] ,\c0|cfg_twr_wire[2] ,\c0|cfg_twr_wire[1] ,\c0|cfg_twr_wire[0] }),
	.afi_mem_clk_disable({\c0|afi_mem_clk_disable[0] }),
	.cfg_dramconfig({cfg_dramconfig_unconnected_wire_23,cfg_dramconfig_unconnected_wire_22,cfg_dramconfig_unconnected_wire_21,\c0|cfg_dramconfig_wire[20] ,\c0|cfg_dramconfig_wire[19] ,\c0|cfg_dramconfig_wire[18] ,\c0|cfg_dramconfig_wire[17] ,\c0|cfg_dramconfig_wire[16] ,
\c0|cfg_dramconfig_wire[15] ,\c0|cfg_dramconfig_wire[14] ,\c0|cfg_dramconfig_wire[13] ,\c0|cfg_dramconfig_wire[12] ,\c0|cfg_dramconfig_wire[11] ,\c0|cfg_dramconfig_wire[10] ,\c0|cfg_dramconfig_wire[9] ,\c0|cfg_dramconfig_wire[8] ,\c0|cfg_dramconfig_wire[7] ,
\c0|cfg_dramconfig_wire[6] ,\c0|cfg_dramconfig_wire[5] ,\c0|cfg_dramconfig_wire[4] ,\c0|cfg_dramconfig_wire[3] ,\c0|cfg_dramconfig_wire[2] ,\c0|cfg_dramconfig_wire[1] ,\c0|cfg_dramconfig_wire[0] }),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ));

terminal_qsys_hps_sdram_p0 p0(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(\p0|umemphy|afi_cal_fail ),
	.afi_cal_success(\p0|umemphy|afi_cal_success ),
	.afi_rdata_valid_0(\p0|umemphy|afi_rdata_valid[0] ),
	.ctl_reset_n(\p0|umemphy|ctl_reset_n ),
	.afi_rdata_0(\p0|umemphy|afi_rdata[0] ),
	.afi_rdata_1(\p0|umemphy|afi_rdata[1] ),
	.afi_rdata_2(\p0|umemphy|afi_rdata[2] ),
	.afi_rdata_3(\p0|umemphy|afi_rdata[3] ),
	.afi_rdata_4(\p0|umemphy|afi_rdata[4] ),
	.afi_rdata_5(\p0|umemphy|afi_rdata[5] ),
	.afi_rdata_6(\p0|umemphy|afi_rdata[6] ),
	.afi_rdata_7(\p0|umemphy|afi_rdata[7] ),
	.afi_rdata_8(\p0|umemphy|afi_rdata[8] ),
	.afi_rdata_9(\p0|umemphy|afi_rdata[9] ),
	.afi_rdata_10(\p0|umemphy|afi_rdata[10] ),
	.afi_rdata_11(\p0|umemphy|afi_rdata[11] ),
	.afi_rdata_12(\p0|umemphy|afi_rdata[12] ),
	.afi_rdata_13(\p0|umemphy|afi_rdata[13] ),
	.afi_rdata_14(\p0|umemphy|afi_rdata[14] ),
	.afi_rdata_15(\p0|umemphy|afi_rdata[15] ),
	.afi_rdata_16(\p0|umemphy|afi_rdata[16] ),
	.afi_rdata_17(\p0|umemphy|afi_rdata[17] ),
	.afi_rdata_18(\p0|umemphy|afi_rdata[18] ),
	.afi_rdata_19(\p0|umemphy|afi_rdata[19] ),
	.afi_rdata_20(\p0|umemphy|afi_rdata[20] ),
	.afi_rdata_21(\p0|umemphy|afi_rdata[21] ),
	.afi_rdata_22(\p0|umemphy|afi_rdata[22] ),
	.afi_rdata_23(\p0|umemphy|afi_rdata[23] ),
	.afi_rdata_24(\p0|umemphy|afi_rdata[24] ),
	.afi_rdata_25(\p0|umemphy|afi_rdata[25] ),
	.afi_rdata_26(\p0|umemphy|afi_rdata[26] ),
	.afi_rdata_27(\p0|umemphy|afi_rdata[27] ),
	.afi_rdata_28(\p0|umemphy|afi_rdata[28] ),
	.afi_rdata_29(\p0|umemphy|afi_rdata[29] ),
	.afi_rdata_30(\p0|umemphy|afi_rdata[30] ),
	.afi_rdata_31(\p0|umemphy|afi_rdata[31] ),
	.afi_rdata_32(\p0|umemphy|afi_rdata[32] ),
	.afi_rdata_33(\p0|umemphy|afi_rdata[33] ),
	.afi_rdata_34(\p0|umemphy|afi_rdata[34] ),
	.afi_rdata_35(\p0|umemphy|afi_rdata[35] ),
	.afi_rdata_36(\p0|umemphy|afi_rdata[36] ),
	.afi_rdata_37(\p0|umemphy|afi_rdata[37] ),
	.afi_rdata_38(\p0|umemphy|afi_rdata[38] ),
	.afi_rdata_39(\p0|umemphy|afi_rdata[39] ),
	.afi_rdata_40(\p0|umemphy|afi_rdata[40] ),
	.afi_rdata_41(\p0|umemphy|afi_rdata[41] ),
	.afi_rdata_42(\p0|umemphy|afi_rdata[42] ),
	.afi_rdata_43(\p0|umemphy|afi_rdata[43] ),
	.afi_rdata_44(\p0|umemphy|afi_rdata[44] ),
	.afi_rdata_45(\p0|umemphy|afi_rdata[45] ),
	.afi_rdata_46(\p0|umemphy|afi_rdata[46] ),
	.afi_rdata_47(\p0|umemphy|afi_rdata[47] ),
	.afi_rdata_48(\p0|umemphy|afi_rdata[48] ),
	.afi_rdata_49(\p0|umemphy|afi_rdata[49] ),
	.afi_rdata_50(\p0|umemphy|afi_rdata[50] ),
	.afi_rdata_51(\p0|umemphy|afi_rdata[51] ),
	.afi_rdata_52(\p0|umemphy|afi_rdata[52] ),
	.afi_rdata_53(\p0|umemphy|afi_rdata[53] ),
	.afi_rdata_54(\p0|umemphy|afi_rdata[54] ),
	.afi_rdata_55(\p0|umemphy|afi_rdata[55] ),
	.afi_rdata_56(\p0|umemphy|afi_rdata[56] ),
	.afi_rdata_57(\p0|umemphy|afi_rdata[57] ),
	.afi_rdata_58(\p0|umemphy|afi_rdata[58] ),
	.afi_rdata_59(\p0|umemphy|afi_rdata[59] ),
	.afi_rdata_60(\p0|umemphy|afi_rdata[60] ),
	.afi_rdata_61(\p0|umemphy|afi_rdata[61] ),
	.afi_rdata_62(\p0|umemphy|afi_rdata[62] ),
	.afi_rdata_63(\p0|umemphy|afi_rdata[63] ),
	.afi_rdata_64(\p0|umemphy|afi_rdata[64] ),
	.afi_rdata_65(\p0|umemphy|afi_rdata[65] ),
	.afi_rdata_66(\p0|umemphy|afi_rdata[66] ),
	.afi_rdata_67(\p0|umemphy|afi_rdata[67] ),
	.afi_rdata_68(\p0|umemphy|afi_rdata[68] ),
	.afi_rdata_69(\p0|umemphy|afi_rdata[69] ),
	.afi_rdata_70(\p0|umemphy|afi_rdata[70] ),
	.afi_rdata_71(\p0|umemphy|afi_rdata[71] ),
	.afi_rdata_72(\p0|umemphy|afi_rdata[72] ),
	.afi_rdata_73(\p0|umemphy|afi_rdata[73] ),
	.afi_rdata_74(\p0|umemphy|afi_rdata[74] ),
	.afi_rdata_75(\p0|umemphy|afi_rdata[75] ),
	.afi_rdata_76(\p0|umemphy|afi_rdata[76] ),
	.afi_rdata_77(\p0|umemphy|afi_rdata[77] ),
	.afi_rdata_78(\p0|umemphy|afi_rdata[78] ),
	.afi_rdata_79(\p0|umemphy|afi_rdata[79] ),
	.afi_wlat_0(\p0|umemphy|afi_wlat[0] ),
	.afi_wlat_1(\p0|umemphy|afi_wlat[1] ),
	.afi_wlat_2(\p0|umemphy|afi_wlat[2] ),
	.afi_wlat_3(\p0|umemphy|afi_wlat[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n_0(\c0|afi_cas_n[0] ),
	.afi_ras_n_0(\c0|afi_ras_n[0] ),
	.afi_rst_n_0(\c0|afi_rst_n[0] ),
	.afi_we_n_0(\c0|afi_we_n[0] ),
	.afi_addr_0(\c0|afi_addr[0] ),
	.afi_addr_1(\c0|afi_addr[1] ),
	.afi_addr_2(\c0|afi_addr[2] ),
	.afi_addr_3(\c0|afi_addr[3] ),
	.afi_addr_4(\c0|afi_addr[4] ),
	.afi_addr_5(\c0|afi_addr[5] ),
	.afi_addr_6(\c0|afi_addr[6] ),
	.afi_addr_7(\c0|afi_addr[7] ),
	.afi_addr_8(\c0|afi_addr[8] ),
	.afi_addr_9(\c0|afi_addr[9] ),
	.afi_addr_10(\c0|afi_addr[10] ),
	.afi_addr_11(\c0|afi_addr[11] ),
	.afi_addr_12(\c0|afi_addr[12] ),
	.afi_addr_13(\c0|afi_addr[13] ),
	.afi_addr_14(\c0|afi_addr[14] ),
	.afi_addr_15(\c0|afi_addr[15] ),
	.afi_addr_16(\c0|afi_addr[16] ),
	.afi_addr_17(\c0|afi_addr[17] ),
	.afi_addr_18(\c0|afi_addr[18] ),
	.afi_addr_19(\c0|afi_addr[19] ),
	.afi_ba_0(\c0|afi_ba[0] ),
	.afi_ba_1(\c0|afi_ba[1] ),
	.afi_ba_2(\c0|afi_ba[2] ),
	.afi_cke_0(\c0|afi_cke[0] ),
	.afi_cke_1(\c0|afi_cke[1] ),
	.afi_cs_n_0(\c0|afi_cs_n[0] ),
	.afi_cs_n_1(\c0|afi_cs_n[1] ),
	.afi_dm_int_0(\c0|afi_dm_int[0] ),
	.afi_dm_int_1(\c0|afi_dm_int[1] ),
	.afi_dm_int_2(\c0|afi_dm_int[2] ),
	.afi_dm_int_3(\c0|afi_dm_int[3] ),
	.afi_dm_int_4(\c0|afi_dm_int[4] ),
	.afi_dm_int_5(\c0|afi_dm_int[5] ),
	.afi_dm_int_6(\c0|afi_dm_int[6] ),
	.afi_dm_int_7(\c0|afi_dm_int[7] ),
	.afi_dm_int_8(\c0|afi_dm_int[8] ),
	.afi_dm_int_9(\c0|afi_dm_int[9] ),
	.afi_dqs_burst_0(\c0|afi_dqs_burst[0] ),
	.afi_dqs_burst_1(\c0|afi_dqs_burst[1] ),
	.afi_dqs_burst_2(\c0|afi_dqs_burst[2] ),
	.afi_dqs_burst_3(\c0|afi_dqs_burst[3] ),
	.afi_dqs_burst_4(\c0|afi_dqs_burst[4] ),
	.afi_odt_0(\c0|afi_odt[0] ),
	.afi_odt_1(\c0|afi_odt[1] ),
	.afi_rdata_en_0(\c0|afi_rdata_en[0] ),
	.afi_rdata_en_1(\c0|afi_rdata_en[1] ),
	.afi_rdata_en_2(\c0|afi_rdata_en[2] ),
	.afi_rdata_en_3(\c0|afi_rdata_en[3] ),
	.afi_rdata_en_4(\c0|afi_rdata_en[4] ),
	.afi_rdata_en_full_0(\c0|afi_rdata_en_full[0] ),
	.afi_rdata_en_full_1(\c0|afi_rdata_en_full[1] ),
	.afi_rdata_en_full_2(\c0|afi_rdata_en_full[2] ),
	.afi_rdata_en_full_3(\c0|afi_rdata_en_full[3] ),
	.afi_rdata_en_full_4(\c0|afi_rdata_en_full[4] ),
	.afi_wdata_int_0(\c0|afi_wdata_int[0] ),
	.afi_wdata_int_1(\c0|afi_wdata_int[1] ),
	.afi_wdata_int_2(\c0|afi_wdata_int[2] ),
	.afi_wdata_int_3(\c0|afi_wdata_int[3] ),
	.afi_wdata_int_4(\c0|afi_wdata_int[4] ),
	.afi_wdata_int_5(\c0|afi_wdata_int[5] ),
	.afi_wdata_int_6(\c0|afi_wdata_int[6] ),
	.afi_wdata_int_7(\c0|afi_wdata_int[7] ),
	.afi_wdata_int_8(\c0|afi_wdata_int[8] ),
	.afi_wdata_int_9(\c0|afi_wdata_int[9] ),
	.afi_wdata_int_10(\c0|afi_wdata_int[10] ),
	.afi_wdata_int_11(\c0|afi_wdata_int[11] ),
	.afi_wdata_int_12(\c0|afi_wdata_int[12] ),
	.afi_wdata_int_13(\c0|afi_wdata_int[13] ),
	.afi_wdata_int_14(\c0|afi_wdata_int[14] ),
	.afi_wdata_int_15(\c0|afi_wdata_int[15] ),
	.afi_wdata_int_16(\c0|afi_wdata_int[16] ),
	.afi_wdata_int_17(\c0|afi_wdata_int[17] ),
	.afi_wdata_int_18(\c0|afi_wdata_int[18] ),
	.afi_wdata_int_19(\c0|afi_wdata_int[19] ),
	.afi_wdata_int_20(\c0|afi_wdata_int[20] ),
	.afi_wdata_int_21(\c0|afi_wdata_int[21] ),
	.afi_wdata_int_22(\c0|afi_wdata_int[22] ),
	.afi_wdata_int_23(\c0|afi_wdata_int[23] ),
	.afi_wdata_int_24(\c0|afi_wdata_int[24] ),
	.afi_wdata_int_25(\c0|afi_wdata_int[25] ),
	.afi_wdata_int_26(\c0|afi_wdata_int[26] ),
	.afi_wdata_int_27(\c0|afi_wdata_int[27] ),
	.afi_wdata_int_28(\c0|afi_wdata_int[28] ),
	.afi_wdata_int_29(\c0|afi_wdata_int[29] ),
	.afi_wdata_int_30(\c0|afi_wdata_int[30] ),
	.afi_wdata_int_31(\c0|afi_wdata_int[31] ),
	.afi_wdata_int_32(\c0|afi_wdata_int[32] ),
	.afi_wdata_int_33(\c0|afi_wdata_int[33] ),
	.afi_wdata_int_34(\c0|afi_wdata_int[34] ),
	.afi_wdata_int_35(\c0|afi_wdata_int[35] ),
	.afi_wdata_int_36(\c0|afi_wdata_int[36] ),
	.afi_wdata_int_37(\c0|afi_wdata_int[37] ),
	.afi_wdata_int_38(\c0|afi_wdata_int[38] ),
	.afi_wdata_int_39(\c0|afi_wdata_int[39] ),
	.afi_wdata_int_40(\c0|afi_wdata_int[40] ),
	.afi_wdata_int_41(\c0|afi_wdata_int[41] ),
	.afi_wdata_int_42(\c0|afi_wdata_int[42] ),
	.afi_wdata_int_43(\c0|afi_wdata_int[43] ),
	.afi_wdata_int_44(\c0|afi_wdata_int[44] ),
	.afi_wdata_int_45(\c0|afi_wdata_int[45] ),
	.afi_wdata_int_46(\c0|afi_wdata_int[46] ),
	.afi_wdata_int_47(\c0|afi_wdata_int[47] ),
	.afi_wdata_int_48(\c0|afi_wdata_int[48] ),
	.afi_wdata_int_49(\c0|afi_wdata_int[49] ),
	.afi_wdata_int_50(\c0|afi_wdata_int[50] ),
	.afi_wdata_int_51(\c0|afi_wdata_int[51] ),
	.afi_wdata_int_52(\c0|afi_wdata_int[52] ),
	.afi_wdata_int_53(\c0|afi_wdata_int[53] ),
	.afi_wdata_int_54(\c0|afi_wdata_int[54] ),
	.afi_wdata_int_55(\c0|afi_wdata_int[55] ),
	.afi_wdata_int_56(\c0|afi_wdata_int[56] ),
	.afi_wdata_int_57(\c0|afi_wdata_int[57] ),
	.afi_wdata_int_58(\c0|afi_wdata_int[58] ),
	.afi_wdata_int_59(\c0|afi_wdata_int[59] ),
	.afi_wdata_int_60(\c0|afi_wdata_int[60] ),
	.afi_wdata_int_61(\c0|afi_wdata_int[61] ),
	.afi_wdata_int_62(\c0|afi_wdata_int[62] ),
	.afi_wdata_int_63(\c0|afi_wdata_int[63] ),
	.afi_wdata_int_64(\c0|afi_wdata_int[64] ),
	.afi_wdata_int_65(\c0|afi_wdata_int[65] ),
	.afi_wdata_int_66(\c0|afi_wdata_int[66] ),
	.afi_wdata_int_67(\c0|afi_wdata_int[67] ),
	.afi_wdata_int_68(\c0|afi_wdata_int[68] ),
	.afi_wdata_int_69(\c0|afi_wdata_int[69] ),
	.afi_wdata_int_70(\c0|afi_wdata_int[70] ),
	.afi_wdata_int_71(\c0|afi_wdata_int[71] ),
	.afi_wdata_int_72(\c0|afi_wdata_int[72] ),
	.afi_wdata_int_73(\c0|afi_wdata_int[73] ),
	.afi_wdata_int_74(\c0|afi_wdata_int[74] ),
	.afi_wdata_int_75(\c0|afi_wdata_int[75] ),
	.afi_wdata_int_76(\c0|afi_wdata_int[76] ),
	.afi_wdata_int_77(\c0|afi_wdata_int[77] ),
	.afi_wdata_int_78(\c0|afi_wdata_int[78] ),
	.afi_wdata_int_79(\c0|afi_wdata_int[79] ),
	.afi_wdata_valid_0(\c0|afi_wdata_valid[0] ),
	.afi_wdata_valid_1(\c0|afi_wdata_valid[1] ),
	.afi_wdata_valid_2(\c0|afi_wdata_valid[2] ),
	.afi_wdata_valid_3(\c0|afi_wdata_valid[3] ),
	.afi_wdata_valid_4(\c0|afi_wdata_valid[4] ),
	.cfg_addlat_wire_0(\c0|cfg_addlat_wire[0] ),
	.cfg_addlat_wire_1(\c0|cfg_addlat_wire[1] ),
	.cfg_addlat_wire_2(\c0|cfg_addlat_wire[2] ),
	.cfg_addlat_wire_3(\c0|cfg_addlat_wire[3] ),
	.cfg_addlat_wire_4(\c0|cfg_addlat_wire[4] ),
	.cfg_bankaddrwidth_wire_0(\c0|cfg_bankaddrwidth_wire[0] ),
	.cfg_bankaddrwidth_wire_1(\c0|cfg_bankaddrwidth_wire[1] ),
	.cfg_bankaddrwidth_wire_2(\c0|cfg_bankaddrwidth_wire[2] ),
	.cfg_caswrlat_wire_0(\c0|cfg_caswrlat_wire[0] ),
	.cfg_caswrlat_wire_1(\c0|cfg_caswrlat_wire[1] ),
	.cfg_caswrlat_wire_2(\c0|cfg_caswrlat_wire[2] ),
	.cfg_caswrlat_wire_3(\c0|cfg_caswrlat_wire[3] ),
	.cfg_coladdrwidth_wire_0(\c0|cfg_coladdrwidth_wire[0] ),
	.cfg_coladdrwidth_wire_1(\c0|cfg_coladdrwidth_wire[1] ),
	.cfg_coladdrwidth_wire_2(\c0|cfg_coladdrwidth_wire[2] ),
	.cfg_coladdrwidth_wire_3(\c0|cfg_coladdrwidth_wire[3] ),
	.cfg_coladdrwidth_wire_4(\c0|cfg_coladdrwidth_wire[4] ),
	.cfg_csaddrwidth_wire_0(\c0|cfg_csaddrwidth_wire[0] ),
	.cfg_csaddrwidth_wire_1(\c0|cfg_csaddrwidth_wire[1] ),
	.cfg_csaddrwidth_wire_2(\c0|cfg_csaddrwidth_wire[2] ),
	.cfg_devicewidth_wire_0(\c0|cfg_devicewidth_wire[0] ),
	.cfg_devicewidth_wire_1(\c0|cfg_devicewidth_wire[1] ),
	.cfg_devicewidth_wire_2(\c0|cfg_devicewidth_wire[2] ),
	.cfg_devicewidth_wire_3(\c0|cfg_devicewidth_wire[3] ),
	.cfg_interfacewidth_wire_0(\c0|cfg_interfacewidth_wire[0] ),
	.cfg_interfacewidth_wire_1(\c0|cfg_interfacewidth_wire[1] ),
	.cfg_interfacewidth_wire_2(\c0|cfg_interfacewidth_wire[2] ),
	.cfg_interfacewidth_wire_3(\c0|cfg_interfacewidth_wire[3] ),
	.cfg_interfacewidth_wire_4(\c0|cfg_interfacewidth_wire[4] ),
	.cfg_interfacewidth_wire_5(\c0|cfg_interfacewidth_wire[5] ),
	.cfg_interfacewidth_wire_6(\c0|cfg_interfacewidth_wire[6] ),
	.cfg_interfacewidth_wire_7(\c0|cfg_interfacewidth_wire[7] ),
	.cfg_rowaddrwidth_wire_0(\c0|cfg_rowaddrwidth_wire[0] ),
	.cfg_rowaddrwidth_wire_1(\c0|cfg_rowaddrwidth_wire[1] ),
	.cfg_rowaddrwidth_wire_2(\c0|cfg_rowaddrwidth_wire[2] ),
	.cfg_rowaddrwidth_wire_3(\c0|cfg_rowaddrwidth_wire[3] ),
	.cfg_rowaddrwidth_wire_4(\c0|cfg_rowaddrwidth_wire[4] ),
	.cfg_tcl_wire_0(\c0|cfg_tcl_wire[0] ),
	.cfg_tcl_wire_1(\c0|cfg_tcl_wire[1] ),
	.cfg_tcl_wire_2(\c0|cfg_tcl_wire[2] ),
	.cfg_tcl_wire_3(\c0|cfg_tcl_wire[3] ),
	.cfg_tcl_wire_4(\c0|cfg_tcl_wire[4] ),
	.cfg_tmrd_wire_0(\c0|cfg_tmrd_wire[0] ),
	.cfg_tmrd_wire_1(\c0|cfg_tmrd_wire[1] ),
	.cfg_tmrd_wire_2(\c0|cfg_tmrd_wire[2] ),
	.cfg_tmrd_wire_3(\c0|cfg_tmrd_wire[3] ),
	.cfg_trefi_wire_0(\c0|cfg_trefi_wire[0] ),
	.cfg_trefi_wire_1(\c0|cfg_trefi_wire[1] ),
	.cfg_trefi_wire_2(\c0|cfg_trefi_wire[2] ),
	.cfg_trefi_wire_3(\c0|cfg_trefi_wire[3] ),
	.cfg_trefi_wire_4(\c0|cfg_trefi_wire[4] ),
	.cfg_trefi_wire_5(\c0|cfg_trefi_wire[5] ),
	.cfg_trefi_wire_6(\c0|cfg_trefi_wire[6] ),
	.cfg_trefi_wire_7(\c0|cfg_trefi_wire[7] ),
	.cfg_trefi_wire_8(\c0|cfg_trefi_wire[8] ),
	.cfg_trefi_wire_9(\c0|cfg_trefi_wire[9] ),
	.cfg_trefi_wire_10(\c0|cfg_trefi_wire[10] ),
	.cfg_trefi_wire_11(\c0|cfg_trefi_wire[11] ),
	.cfg_trefi_wire_12(\c0|cfg_trefi_wire[12] ),
	.cfg_trfc_wire_0(\c0|cfg_trfc_wire[0] ),
	.cfg_trfc_wire_1(\c0|cfg_trfc_wire[1] ),
	.cfg_trfc_wire_2(\c0|cfg_trfc_wire[2] ),
	.cfg_trfc_wire_3(\c0|cfg_trfc_wire[3] ),
	.cfg_trfc_wire_4(\c0|cfg_trfc_wire[4] ),
	.cfg_trfc_wire_5(\c0|cfg_trfc_wire[5] ),
	.cfg_trfc_wire_6(\c0|cfg_trfc_wire[6] ),
	.cfg_trfc_wire_7(\c0|cfg_trfc_wire[7] ),
	.cfg_twr_wire_0(\c0|cfg_twr_wire[0] ),
	.cfg_twr_wire_1(\c0|cfg_twr_wire[1] ),
	.cfg_twr_wire_2(\c0|cfg_twr_wire[2] ),
	.cfg_twr_wire_3(\c0|cfg_twr_wire[3] ),
	.afi_mem_clk_disable_0(\c0|afi_mem_clk_disable[0] ),
	.cfg_dramconfig_wire_0(\c0|cfg_dramconfig_wire[0] ),
	.cfg_dramconfig_wire_1(\c0|cfg_dramconfig_wire[1] ),
	.cfg_dramconfig_wire_2(\c0|cfg_dramconfig_wire[2] ),
	.cfg_dramconfig_wire_3(\c0|cfg_dramconfig_wire[3] ),
	.cfg_dramconfig_wire_4(\c0|cfg_dramconfig_wire[4] ),
	.cfg_dramconfig_wire_5(\c0|cfg_dramconfig_wire[5] ),
	.cfg_dramconfig_wire_6(\c0|cfg_dramconfig_wire[6] ),
	.cfg_dramconfig_wire_7(\c0|cfg_dramconfig_wire[7] ),
	.cfg_dramconfig_wire_8(\c0|cfg_dramconfig_wire[8] ),
	.cfg_dramconfig_wire_9(\c0|cfg_dramconfig_wire[9] ),
	.cfg_dramconfig_wire_10(\c0|cfg_dramconfig_wire[10] ),
	.cfg_dramconfig_wire_11(\c0|cfg_dramconfig_wire[11] ),
	.cfg_dramconfig_wire_12(\c0|cfg_dramconfig_wire[12] ),
	.cfg_dramconfig_wire_13(\c0|cfg_dramconfig_wire[13] ),
	.cfg_dramconfig_wire_14(\c0|cfg_dramconfig_wire[14] ),
	.cfg_dramconfig_wire_15(\c0|cfg_dramconfig_wire[15] ),
	.cfg_dramconfig_wire_16(\c0|cfg_dramconfig_wire[16] ),
	.cfg_dramconfig_wire_17(\c0|cfg_dramconfig_wire[17] ),
	.cfg_dramconfig_wire_18(\c0|cfg_dramconfig_wire[18] ),
	.cfg_dramconfig_wire_19(\c0|cfg_dramconfig_wire[19] ),
	.cfg_dramconfig_wire_20(\c0|cfg_dramconfig_wire[20] ),
	.ctl_clk(\p0|umemphy|memphy_ldc|leveled_dqs_clocks[0] ),
	.dll_delayctrl_0(\dll|dll_delayctrl[0] ),
	.dll_delayctrl_1(\dll|dll_delayctrl[1] ),
	.dll_delayctrl_2(\dll|dll_delayctrl[2] ),
	.dll_delayctrl_3(\dll|dll_delayctrl[3] ),
	.dll_delayctrl_4(\dll|dll_delayctrl[4] ),
	.dll_delayctrl_5(\dll|dll_delayctrl[5] ),
	.dll_delayctrl_6(\dll|dll_delayctrl[6] ),
	.GND_port(GND_port));

terminal_qsys_hps_sdram_pll pll(
	.pll_mem_clk(\pll|afi_clk ),
	.pll_write_clk(\pll|pll_write_clk ));

endmodule

module terminal_qsys_altera_mem_if_dll_cyclonev (
	clk,
	dll_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	[6:0] dll_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [6:0] dll_wys_m_DELAYCTRLOUT_bus;

assign dll_delayctrl[0] = dll_wys_m_DELAYCTRLOUT_bus[0];
assign dll_delayctrl[1] = dll_wys_m_DELAYCTRLOUT_bus[1];
assign dll_delayctrl[2] = dll_wys_m_DELAYCTRLOUT_bus[2];
assign dll_delayctrl[3] = dll_wys_m_DELAYCTRLOUT_bus[3];
assign dll_delayctrl[4] = dll_wys_m_DELAYCTRLOUT_bus[4];
assign dll_delayctrl[5] = dll_wys_m_DELAYCTRLOUT_bus[5];
assign dll_delayctrl[6] = dll_wys_m_DELAYCTRLOUT_bus[6];

cyclonev_dll dll_wys_m(
	.clk(clk),
	.aload(vcc),
	.upndnin(gnd),
	.upndninclkena(gnd),
	.dqsupdate(),
	.upndnout(),
	.delayctrlout(dll_wys_m_DELAYCTRLOUT_bus));
defparam dll_wys_m.delayctrlout_mode = "normal";
defparam dll_wys_m.input_frequency = "2500 ps";
defparam dll_wys_m.jitter_reduction = "true";
defparam dll_wys_m.sim_buffer_delay_increment = 10;
defparam dll_wys_m.sim_buffer_intrinsic_delay = 175;
defparam dll_wys_m.sim_valid_lock = 16;
defparam dll_wys_m.sim_valid_lockcount = 0;
defparam dll_wys_m.static_delay_ctrl = 8;
defparam dll_wys_m.upndnout_mode = "clock";
defparam dll_wys_m.use_upndnin = "false";
defparam dll_wys_m.use_upndninclkena = "false";

endmodule

module terminal_qsys_altera_mem_if_hard_memory_controller_top_cyclonev (
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk)/* synthesis synthesis_greybox=0 */;
input 	afi_cal_fail;
input 	afi_cal_success;
input 	[0:0] afi_rdata_valid;
input 	ctl_reset_n;
input 	[79:0] afi_rdata;
input 	[3:0] afi_wlat;
output 	[0:0] afi_cas_n;
output 	[0:0] afi_ras_n;
output 	[0:0] afi_rst_n;
output 	[0:0] afi_we_n;
output 	[19:0] afi_addr;
output 	[2:0] afi_ba;
output 	[1:0] afi_cke;
output 	[1:0] afi_cs_n;
output 	[9:0] afi_dm;
output 	[4:0] afi_dqs_burst;
output 	[1:0] afi_odt;
output 	[4:0] afi_rdata_en;
output 	[4:0] afi_rdata_en_full;
output 	[79:0] afi_wdata;
output 	[4:0] afi_wdata_valid;
output 	[7:0] cfg_addlat;
output 	[7:0] cfg_bankaddrwidth;
output 	[7:0] cfg_caswrlat;
output 	[7:0] cfg_coladdrwidth;
output 	[7:0] cfg_csaddrwidth;
output 	[7:0] cfg_devicewidth;
output 	[7:0] cfg_interfacewidth;
output 	[7:0] cfg_rowaddrwidth;
output 	[7:0] cfg_tcl;
output 	[7:0] cfg_tmrd;
output 	[15:0] cfg_trefi;
output 	[7:0] cfg_trfc;
output 	[7:0] cfg_twr;
output 	[0:0] afi_mem_clk_disable;
output 	[23:0] cfg_dramconfig;
input 	ctl_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [19:0] hmc_inst_AFIADDR_bus;
wire [2:0] hmc_inst_AFIBA_bus;
wire [1:0] hmc_inst_AFICKE_bus;
wire [1:0] hmc_inst_AFICSN_bus;
wire [9:0] hmc_inst_AFIDM_bus;
wire [4:0] hmc_inst_AFIDQSBURST_bus;
wire [1:0] hmc_inst_AFIODT_bus;
wire [4:0] hmc_inst_AFIRDATAEN_bus;
wire [4:0] hmc_inst_AFIRDATAENFULL_bus;
wire [79:0] hmc_inst_AFIWDATA_bus;
wire [4:0] hmc_inst_AFIWDATAVALID_bus;
wire [4:0] hmc_inst_CFGADDLAT_bus;
wire [2:0] hmc_inst_CFGBANKADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGCASWRLAT_bus;
wire [4:0] hmc_inst_CFGCOLADDRWIDTH_bus;
wire [2:0] hmc_inst_CFGCSADDRWIDTH_bus;
wire [3:0] hmc_inst_CFGDEVICEWIDTH_bus;
wire [7:0] hmc_inst_CFGINTERFACEWIDTH_bus;
wire [4:0] hmc_inst_CFGROWADDRWIDTH_bus;
wire [4:0] hmc_inst_CFGTCL_bus;
wire [3:0] hmc_inst_CFGTMRD_bus;
wire [12:0] hmc_inst_CFGTREFI_bus;
wire [7:0] hmc_inst_CFGTRFC_bus;
wire [3:0] hmc_inst_CFGTWR_bus;
wire [1:0] hmc_inst_CTLMEMCLKDISABLE_bus;
wire [20:0] hmc_inst_DRAMCONFIG_bus;

assign afi_addr[0] = hmc_inst_AFIADDR_bus[0];
assign afi_addr[1] = hmc_inst_AFIADDR_bus[1];
assign afi_addr[2] = hmc_inst_AFIADDR_bus[2];
assign afi_addr[3] = hmc_inst_AFIADDR_bus[3];
assign afi_addr[4] = hmc_inst_AFIADDR_bus[4];
assign afi_addr[5] = hmc_inst_AFIADDR_bus[5];
assign afi_addr[6] = hmc_inst_AFIADDR_bus[6];
assign afi_addr[7] = hmc_inst_AFIADDR_bus[7];
assign afi_addr[8] = hmc_inst_AFIADDR_bus[8];
assign afi_addr[9] = hmc_inst_AFIADDR_bus[9];
assign afi_addr[10] = hmc_inst_AFIADDR_bus[10];
assign afi_addr[11] = hmc_inst_AFIADDR_bus[11];
assign afi_addr[12] = hmc_inst_AFIADDR_bus[12];
assign afi_addr[13] = hmc_inst_AFIADDR_bus[13];
assign afi_addr[14] = hmc_inst_AFIADDR_bus[14];
assign afi_addr[15] = hmc_inst_AFIADDR_bus[15];
assign afi_addr[16] = hmc_inst_AFIADDR_bus[16];
assign afi_addr[17] = hmc_inst_AFIADDR_bus[17];
assign afi_addr[18] = hmc_inst_AFIADDR_bus[18];
assign afi_addr[19] = hmc_inst_AFIADDR_bus[19];

assign afi_ba[0] = hmc_inst_AFIBA_bus[0];
assign afi_ba[1] = hmc_inst_AFIBA_bus[1];
assign afi_ba[2] = hmc_inst_AFIBA_bus[2];

assign afi_cke[0] = hmc_inst_AFICKE_bus[0];
assign afi_cke[1] = hmc_inst_AFICKE_bus[1];

assign afi_cs_n[0] = hmc_inst_AFICSN_bus[0];
assign afi_cs_n[1] = hmc_inst_AFICSN_bus[1];

assign afi_dm[0] = hmc_inst_AFIDM_bus[0];
assign afi_dm[1] = hmc_inst_AFIDM_bus[1];
assign afi_dm[2] = hmc_inst_AFIDM_bus[2];
assign afi_dm[3] = hmc_inst_AFIDM_bus[3];
assign afi_dm[4] = hmc_inst_AFIDM_bus[4];
assign afi_dm[5] = hmc_inst_AFIDM_bus[5];
assign afi_dm[6] = hmc_inst_AFIDM_bus[6];
assign afi_dm[7] = hmc_inst_AFIDM_bus[7];
assign afi_dm[8] = hmc_inst_AFIDM_bus[8];
assign afi_dm[9] = hmc_inst_AFIDM_bus[9];

assign afi_dqs_burst[0] = hmc_inst_AFIDQSBURST_bus[0];
assign afi_dqs_burst[1] = hmc_inst_AFIDQSBURST_bus[1];
assign afi_dqs_burst[2] = hmc_inst_AFIDQSBURST_bus[2];
assign afi_dqs_burst[3] = hmc_inst_AFIDQSBURST_bus[3];
assign afi_dqs_burst[4] = hmc_inst_AFIDQSBURST_bus[4];

assign afi_odt[0] = hmc_inst_AFIODT_bus[0];
assign afi_odt[1] = hmc_inst_AFIODT_bus[1];

assign afi_rdata_en[0] = hmc_inst_AFIRDATAEN_bus[0];
assign afi_rdata_en[1] = hmc_inst_AFIRDATAEN_bus[1];
assign afi_rdata_en[2] = hmc_inst_AFIRDATAEN_bus[2];
assign afi_rdata_en[3] = hmc_inst_AFIRDATAEN_bus[3];
assign afi_rdata_en[4] = hmc_inst_AFIRDATAEN_bus[4];

assign afi_rdata_en_full[0] = hmc_inst_AFIRDATAENFULL_bus[0];
assign afi_rdata_en_full[1] = hmc_inst_AFIRDATAENFULL_bus[1];
assign afi_rdata_en_full[2] = hmc_inst_AFIRDATAENFULL_bus[2];
assign afi_rdata_en_full[3] = hmc_inst_AFIRDATAENFULL_bus[3];
assign afi_rdata_en_full[4] = hmc_inst_AFIRDATAENFULL_bus[4];

assign afi_wdata[0] = hmc_inst_AFIWDATA_bus[0];
assign afi_wdata[1] = hmc_inst_AFIWDATA_bus[1];
assign afi_wdata[2] = hmc_inst_AFIWDATA_bus[2];
assign afi_wdata[3] = hmc_inst_AFIWDATA_bus[3];
assign afi_wdata[4] = hmc_inst_AFIWDATA_bus[4];
assign afi_wdata[5] = hmc_inst_AFIWDATA_bus[5];
assign afi_wdata[6] = hmc_inst_AFIWDATA_bus[6];
assign afi_wdata[7] = hmc_inst_AFIWDATA_bus[7];
assign afi_wdata[8] = hmc_inst_AFIWDATA_bus[8];
assign afi_wdata[9] = hmc_inst_AFIWDATA_bus[9];
assign afi_wdata[10] = hmc_inst_AFIWDATA_bus[10];
assign afi_wdata[11] = hmc_inst_AFIWDATA_bus[11];
assign afi_wdata[12] = hmc_inst_AFIWDATA_bus[12];
assign afi_wdata[13] = hmc_inst_AFIWDATA_bus[13];
assign afi_wdata[14] = hmc_inst_AFIWDATA_bus[14];
assign afi_wdata[15] = hmc_inst_AFIWDATA_bus[15];
assign afi_wdata[16] = hmc_inst_AFIWDATA_bus[16];
assign afi_wdata[17] = hmc_inst_AFIWDATA_bus[17];
assign afi_wdata[18] = hmc_inst_AFIWDATA_bus[18];
assign afi_wdata[19] = hmc_inst_AFIWDATA_bus[19];
assign afi_wdata[20] = hmc_inst_AFIWDATA_bus[20];
assign afi_wdata[21] = hmc_inst_AFIWDATA_bus[21];
assign afi_wdata[22] = hmc_inst_AFIWDATA_bus[22];
assign afi_wdata[23] = hmc_inst_AFIWDATA_bus[23];
assign afi_wdata[24] = hmc_inst_AFIWDATA_bus[24];
assign afi_wdata[25] = hmc_inst_AFIWDATA_bus[25];
assign afi_wdata[26] = hmc_inst_AFIWDATA_bus[26];
assign afi_wdata[27] = hmc_inst_AFIWDATA_bus[27];
assign afi_wdata[28] = hmc_inst_AFIWDATA_bus[28];
assign afi_wdata[29] = hmc_inst_AFIWDATA_bus[29];
assign afi_wdata[30] = hmc_inst_AFIWDATA_bus[30];
assign afi_wdata[31] = hmc_inst_AFIWDATA_bus[31];
assign afi_wdata[32] = hmc_inst_AFIWDATA_bus[32];
assign afi_wdata[33] = hmc_inst_AFIWDATA_bus[33];
assign afi_wdata[34] = hmc_inst_AFIWDATA_bus[34];
assign afi_wdata[35] = hmc_inst_AFIWDATA_bus[35];
assign afi_wdata[36] = hmc_inst_AFIWDATA_bus[36];
assign afi_wdata[37] = hmc_inst_AFIWDATA_bus[37];
assign afi_wdata[38] = hmc_inst_AFIWDATA_bus[38];
assign afi_wdata[39] = hmc_inst_AFIWDATA_bus[39];
assign afi_wdata[40] = hmc_inst_AFIWDATA_bus[40];
assign afi_wdata[41] = hmc_inst_AFIWDATA_bus[41];
assign afi_wdata[42] = hmc_inst_AFIWDATA_bus[42];
assign afi_wdata[43] = hmc_inst_AFIWDATA_bus[43];
assign afi_wdata[44] = hmc_inst_AFIWDATA_bus[44];
assign afi_wdata[45] = hmc_inst_AFIWDATA_bus[45];
assign afi_wdata[46] = hmc_inst_AFIWDATA_bus[46];
assign afi_wdata[47] = hmc_inst_AFIWDATA_bus[47];
assign afi_wdata[48] = hmc_inst_AFIWDATA_bus[48];
assign afi_wdata[49] = hmc_inst_AFIWDATA_bus[49];
assign afi_wdata[50] = hmc_inst_AFIWDATA_bus[50];
assign afi_wdata[51] = hmc_inst_AFIWDATA_bus[51];
assign afi_wdata[52] = hmc_inst_AFIWDATA_bus[52];
assign afi_wdata[53] = hmc_inst_AFIWDATA_bus[53];
assign afi_wdata[54] = hmc_inst_AFIWDATA_bus[54];
assign afi_wdata[55] = hmc_inst_AFIWDATA_bus[55];
assign afi_wdata[56] = hmc_inst_AFIWDATA_bus[56];
assign afi_wdata[57] = hmc_inst_AFIWDATA_bus[57];
assign afi_wdata[58] = hmc_inst_AFIWDATA_bus[58];
assign afi_wdata[59] = hmc_inst_AFIWDATA_bus[59];
assign afi_wdata[60] = hmc_inst_AFIWDATA_bus[60];
assign afi_wdata[61] = hmc_inst_AFIWDATA_bus[61];
assign afi_wdata[62] = hmc_inst_AFIWDATA_bus[62];
assign afi_wdata[63] = hmc_inst_AFIWDATA_bus[63];
assign afi_wdata[64] = hmc_inst_AFIWDATA_bus[64];
assign afi_wdata[65] = hmc_inst_AFIWDATA_bus[65];
assign afi_wdata[66] = hmc_inst_AFIWDATA_bus[66];
assign afi_wdata[67] = hmc_inst_AFIWDATA_bus[67];
assign afi_wdata[68] = hmc_inst_AFIWDATA_bus[68];
assign afi_wdata[69] = hmc_inst_AFIWDATA_bus[69];
assign afi_wdata[70] = hmc_inst_AFIWDATA_bus[70];
assign afi_wdata[71] = hmc_inst_AFIWDATA_bus[71];
assign afi_wdata[72] = hmc_inst_AFIWDATA_bus[72];
assign afi_wdata[73] = hmc_inst_AFIWDATA_bus[73];
assign afi_wdata[74] = hmc_inst_AFIWDATA_bus[74];
assign afi_wdata[75] = hmc_inst_AFIWDATA_bus[75];
assign afi_wdata[76] = hmc_inst_AFIWDATA_bus[76];
assign afi_wdata[77] = hmc_inst_AFIWDATA_bus[77];
assign afi_wdata[78] = hmc_inst_AFIWDATA_bus[78];
assign afi_wdata[79] = hmc_inst_AFIWDATA_bus[79];

assign afi_wdata_valid[0] = hmc_inst_AFIWDATAVALID_bus[0];
assign afi_wdata_valid[1] = hmc_inst_AFIWDATAVALID_bus[1];
assign afi_wdata_valid[2] = hmc_inst_AFIWDATAVALID_bus[2];
assign afi_wdata_valid[3] = hmc_inst_AFIWDATAVALID_bus[3];
assign afi_wdata_valid[4] = hmc_inst_AFIWDATAVALID_bus[4];

assign cfg_addlat[0] = hmc_inst_CFGADDLAT_bus[0];
assign cfg_addlat[1] = hmc_inst_CFGADDLAT_bus[1];
assign cfg_addlat[2] = hmc_inst_CFGADDLAT_bus[2];
assign cfg_addlat[3] = hmc_inst_CFGADDLAT_bus[3];
assign cfg_addlat[4] = hmc_inst_CFGADDLAT_bus[4];

assign cfg_bankaddrwidth[0] = hmc_inst_CFGBANKADDRWIDTH_bus[0];
assign cfg_bankaddrwidth[1] = hmc_inst_CFGBANKADDRWIDTH_bus[1];
assign cfg_bankaddrwidth[2] = hmc_inst_CFGBANKADDRWIDTH_bus[2];

assign cfg_caswrlat[0] = hmc_inst_CFGCASWRLAT_bus[0];
assign cfg_caswrlat[1] = hmc_inst_CFGCASWRLAT_bus[1];
assign cfg_caswrlat[2] = hmc_inst_CFGCASWRLAT_bus[2];
assign cfg_caswrlat[3] = hmc_inst_CFGCASWRLAT_bus[3];

assign cfg_coladdrwidth[0] = hmc_inst_CFGCOLADDRWIDTH_bus[0];
assign cfg_coladdrwidth[1] = hmc_inst_CFGCOLADDRWIDTH_bus[1];
assign cfg_coladdrwidth[2] = hmc_inst_CFGCOLADDRWIDTH_bus[2];
assign cfg_coladdrwidth[3] = hmc_inst_CFGCOLADDRWIDTH_bus[3];
assign cfg_coladdrwidth[4] = hmc_inst_CFGCOLADDRWIDTH_bus[4];

assign cfg_csaddrwidth[0] = hmc_inst_CFGCSADDRWIDTH_bus[0];
assign cfg_csaddrwidth[1] = hmc_inst_CFGCSADDRWIDTH_bus[1];
assign cfg_csaddrwidth[2] = hmc_inst_CFGCSADDRWIDTH_bus[2];

assign cfg_devicewidth[0] = hmc_inst_CFGDEVICEWIDTH_bus[0];
assign cfg_devicewidth[1] = hmc_inst_CFGDEVICEWIDTH_bus[1];
assign cfg_devicewidth[2] = hmc_inst_CFGDEVICEWIDTH_bus[2];
assign cfg_devicewidth[3] = hmc_inst_CFGDEVICEWIDTH_bus[3];

assign cfg_interfacewidth[0] = hmc_inst_CFGINTERFACEWIDTH_bus[0];
assign cfg_interfacewidth[1] = hmc_inst_CFGINTERFACEWIDTH_bus[1];
assign cfg_interfacewidth[2] = hmc_inst_CFGINTERFACEWIDTH_bus[2];
assign cfg_interfacewidth[3] = hmc_inst_CFGINTERFACEWIDTH_bus[3];
assign cfg_interfacewidth[4] = hmc_inst_CFGINTERFACEWIDTH_bus[4];
assign cfg_interfacewidth[5] = hmc_inst_CFGINTERFACEWIDTH_bus[5];
assign cfg_interfacewidth[6] = hmc_inst_CFGINTERFACEWIDTH_bus[6];
assign cfg_interfacewidth[7] = hmc_inst_CFGINTERFACEWIDTH_bus[7];

assign cfg_rowaddrwidth[0] = hmc_inst_CFGROWADDRWIDTH_bus[0];
assign cfg_rowaddrwidth[1] = hmc_inst_CFGROWADDRWIDTH_bus[1];
assign cfg_rowaddrwidth[2] = hmc_inst_CFGROWADDRWIDTH_bus[2];
assign cfg_rowaddrwidth[3] = hmc_inst_CFGROWADDRWIDTH_bus[3];
assign cfg_rowaddrwidth[4] = hmc_inst_CFGROWADDRWIDTH_bus[4];

assign cfg_tcl[0] = hmc_inst_CFGTCL_bus[0];
assign cfg_tcl[1] = hmc_inst_CFGTCL_bus[1];
assign cfg_tcl[2] = hmc_inst_CFGTCL_bus[2];
assign cfg_tcl[3] = hmc_inst_CFGTCL_bus[3];
assign cfg_tcl[4] = hmc_inst_CFGTCL_bus[4];

assign cfg_tmrd[0] = hmc_inst_CFGTMRD_bus[0];
assign cfg_tmrd[1] = hmc_inst_CFGTMRD_bus[1];
assign cfg_tmrd[2] = hmc_inst_CFGTMRD_bus[2];
assign cfg_tmrd[3] = hmc_inst_CFGTMRD_bus[3];

assign cfg_trefi[0] = hmc_inst_CFGTREFI_bus[0];
assign cfg_trefi[1] = hmc_inst_CFGTREFI_bus[1];
assign cfg_trefi[2] = hmc_inst_CFGTREFI_bus[2];
assign cfg_trefi[3] = hmc_inst_CFGTREFI_bus[3];
assign cfg_trefi[4] = hmc_inst_CFGTREFI_bus[4];
assign cfg_trefi[5] = hmc_inst_CFGTREFI_bus[5];
assign cfg_trefi[6] = hmc_inst_CFGTREFI_bus[6];
assign cfg_trefi[7] = hmc_inst_CFGTREFI_bus[7];
assign cfg_trefi[8] = hmc_inst_CFGTREFI_bus[8];
assign cfg_trefi[9] = hmc_inst_CFGTREFI_bus[9];
assign cfg_trefi[10] = hmc_inst_CFGTREFI_bus[10];
assign cfg_trefi[11] = hmc_inst_CFGTREFI_bus[11];
assign cfg_trefi[12] = hmc_inst_CFGTREFI_bus[12];

assign cfg_trfc[0] = hmc_inst_CFGTRFC_bus[0];
assign cfg_trfc[1] = hmc_inst_CFGTRFC_bus[1];
assign cfg_trfc[2] = hmc_inst_CFGTRFC_bus[2];
assign cfg_trfc[3] = hmc_inst_CFGTRFC_bus[3];
assign cfg_trfc[4] = hmc_inst_CFGTRFC_bus[4];
assign cfg_trfc[5] = hmc_inst_CFGTRFC_bus[5];
assign cfg_trfc[6] = hmc_inst_CFGTRFC_bus[6];
assign cfg_trfc[7] = hmc_inst_CFGTRFC_bus[7];

assign cfg_twr[0] = hmc_inst_CFGTWR_bus[0];
assign cfg_twr[1] = hmc_inst_CFGTWR_bus[1];
assign cfg_twr[2] = hmc_inst_CFGTWR_bus[2];
assign cfg_twr[3] = hmc_inst_CFGTWR_bus[3];

assign afi_mem_clk_disable[0] = hmc_inst_CTLMEMCLKDISABLE_bus[0];

assign cfg_dramconfig[0] = hmc_inst_DRAMCONFIG_bus[0];
assign cfg_dramconfig[1] = hmc_inst_DRAMCONFIG_bus[1];
assign cfg_dramconfig[2] = hmc_inst_DRAMCONFIG_bus[2];
assign cfg_dramconfig[3] = hmc_inst_DRAMCONFIG_bus[3];
assign cfg_dramconfig[4] = hmc_inst_DRAMCONFIG_bus[4];
assign cfg_dramconfig[5] = hmc_inst_DRAMCONFIG_bus[5];
assign cfg_dramconfig[6] = hmc_inst_DRAMCONFIG_bus[6];
assign cfg_dramconfig[7] = hmc_inst_DRAMCONFIG_bus[7];
assign cfg_dramconfig[8] = hmc_inst_DRAMCONFIG_bus[8];
assign cfg_dramconfig[9] = hmc_inst_DRAMCONFIG_bus[9];
assign cfg_dramconfig[10] = hmc_inst_DRAMCONFIG_bus[10];
assign cfg_dramconfig[11] = hmc_inst_DRAMCONFIG_bus[11];
assign cfg_dramconfig[12] = hmc_inst_DRAMCONFIG_bus[12];
assign cfg_dramconfig[13] = hmc_inst_DRAMCONFIG_bus[13];
assign cfg_dramconfig[14] = hmc_inst_DRAMCONFIG_bus[14];
assign cfg_dramconfig[15] = hmc_inst_DRAMCONFIG_bus[15];
assign cfg_dramconfig[16] = hmc_inst_DRAMCONFIG_bus[16];
assign cfg_dramconfig[17] = hmc_inst_DRAMCONFIG_bus[17];
assign cfg_dramconfig[18] = hmc_inst_DRAMCONFIG_bus[18];
assign cfg_dramconfig[19] = hmc_inst_DRAMCONFIG_bus[19];
assign cfg_dramconfig[20] = hmc_inst_DRAMCONFIG_bus[20];

cyclonev_hmc hmc_inst(
	.afirdatavalid(afi_rdata_valid[0]),
	.csrclk(gnd),
	.csrdin(gnd),
	.csren(gnd),
	.ctlcalfail(afi_cal_fail),
	.ctlcalsuccess(afi_cal_success),
	.ctlclk(ctl_clk),
	.ctlresetn(ctl_reset_n),
	.globalresetn(gnd),
	.iavstcmdresetn0(vcc),
	.iavstcmdresetn1(vcc),
	.iavstcmdresetn2(vcc),
	.iavstcmdresetn3(vcc),
	.iavstcmdresetn4(vcc),
	.iavstcmdresetn5(vcc),
	.iavstrdclk0(gnd),
	.iavstrdclk1(gnd),
	.iavstrdclk2(gnd),
	.iavstrdclk3(gnd),
	.iavstrdready0(vcc),
	.iavstrdready1(vcc),
	.iavstrdready2(vcc),
	.iavstrdready3(vcc),
	.iavstrdresetn0(vcc),
	.iavstrdresetn1(vcc),
	.iavstrdresetn2(vcc),
	.iavstrdresetn3(vcc),
	.iavstwrackready0(vcc),
	.iavstwrackready1(vcc),
	.iavstwrackready2(vcc),
	.iavstwrackready3(vcc),
	.iavstwrackready4(vcc),
	.iavstwrackready5(vcc),
	.iavstwrclk0(gnd),
	.iavstwrclk1(gnd),
	.iavstwrclk2(gnd),
	.iavstwrclk3(gnd),
	.iavstwrresetn0(vcc),
	.iavstwrresetn1(vcc),
	.iavstwrresetn2(vcc),
	.iavstwrresetn3(vcc),
	.localdeeppowerdnreq(gnd),
	.localrefreshreq(gnd),
	.localselfrfshreq(gnd),
	.mmrbe(gnd),
	.mmrburstbegin(vcc),
	.mmrclk(gnd),
	.mmrreadreq(gnd),
	.mmrresetn(vcc),
	.mmrwritereq(gnd),
	.portclk0(gnd),
	.portclk1(gnd),
	.portclk2(gnd),
	.portclk3(gnd),
	.portclk4(gnd),
	.portclk5(gnd),
	.scanenable(gnd),
	.scbe(gnd),
	.scburstbegin(gnd),
	.scclk(gnd),
	.screadreq(gnd),
	.scresetn(vcc),
	.scwritereq(gnd),
	.afirdata({afi_rdata[79],afi_rdata[78],afi_rdata[77],afi_rdata[76],afi_rdata[75],afi_rdata[74],afi_rdata[73],afi_rdata[72],afi_rdata[71],afi_rdata[70],afi_rdata[69],afi_rdata[68],afi_rdata[67],afi_rdata[66],afi_rdata[65],afi_rdata[64],afi_rdata[63],afi_rdata[62],afi_rdata[61],afi_rdata[60],afi_rdata[59],afi_rdata[58],afi_rdata[57],afi_rdata[56],afi_rdata[55],afi_rdata[54],afi_rdata[53],afi_rdata[52],
afi_rdata[51],afi_rdata[50],afi_rdata[49],afi_rdata[48],afi_rdata[47],afi_rdata[46],afi_rdata[45],afi_rdata[44],afi_rdata[43],afi_rdata[42],afi_rdata[41],afi_rdata[40],afi_rdata[39],afi_rdata[38],afi_rdata[37],afi_rdata[36],afi_rdata[35],afi_rdata[34],afi_rdata[33],afi_rdata[32],afi_rdata[31],afi_rdata[30],afi_rdata[29],afi_rdata[28],afi_rdata[27],afi_rdata[26],afi_rdata[25],afi_rdata[24],
afi_rdata[23],afi_rdata[22],afi_rdata[21],afi_rdata[20],afi_rdata[19],afi_rdata[18],afi_rdata[17],afi_rdata[16],afi_rdata[15],afi_rdata[14],afi_rdata[13],afi_rdata[12],afi_rdata[11],afi_rdata[10],afi_rdata[9],afi_rdata[8],afi_rdata[7],afi_rdata[6],afi_rdata[5],afi_rdata[4],afi_rdata[3],afi_rdata[2],afi_rdata[1],afi_rdata[0]}),
	.afiseqbusy({gnd,gnd}),
	.afiwlat({afi_wlat[3],afi_wlat[2],afi_wlat[1],afi_wlat[0]}),
	.bondingin1({gnd,gnd,gnd,gnd}),
	.bondingin2({gnd,gnd,gnd,gnd,gnd,gnd}),
	.bondingin3({gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata4({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstcmddata5({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata0({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata1({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata2({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iavstwrdata3({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.localdeeppowerdnchip({gnd,gnd}),
	.localrefreshchip({gnd,gnd}),
	.localselfrfshchip({gnd,gnd}),
	.mmraddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.mmrburstcount({gnd,vcc}),
	.mmrwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.scburstcount({gnd,gnd}),
	.scwdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.aficasn(afi_cas_n[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.csrdout(),
	.ctlcalreq(),
	.ctlinitreq(),
	.localdeeppowerdnack(),
	.localinitdone(),
	.localpowerdownack(),
	.localrefreshack(),
	.localselfrfshack(),
	.localstsctlempty(),
	.mmrrdatavalid(),
	.mmrwaitrequest(),
	.oammready0(),
	.oammready1(),
	.oammready2(),
	.oammready3(),
	.oammready4(),
	.oammready5(),
	.ordavstvalid0(),
	.ordavstvalid1(),
	.ordavstvalid2(),
	.ordavstvalid3(),
	.owrackavstdata0(),
	.owrackavstdata1(),
	.owrackavstdata2(),
	.owrackavstdata3(),
	.owrackavstdata4(),
	.owrackavstdata5(),
	.owrackavstvalid0(),
	.owrackavstvalid1(),
	.owrackavstvalid2(),
	.owrackavstvalid3(),
	.owrackavstvalid4(),
	.owrackavstvalid5(),
	.scrdatavalid(),
	.scwaitrequest(),
	.afiaddr(hmc_inst_AFIADDR_bus),
	.afiba(hmc_inst_AFIBA_bus),
	.aficke(hmc_inst_AFICKE_bus),
	.aficsn(hmc_inst_AFICSN_bus),
	.afictllongidle(),
	.afictlrefreshdone(),
	.afidm(hmc_inst_AFIDM_bus),
	.afidqsburst(hmc_inst_AFIDQSBURST_bus),
	.afiodt(hmc_inst_AFIODT_bus),
	.afirdataen(hmc_inst_AFIRDATAEN_bus),
	.afirdataenfull(hmc_inst_AFIRDATAENFULL_bus),
	.afiwdata(hmc_inst_AFIWDATA_bus),
	.afiwdatavalid(hmc_inst_AFIWDATAVALID_bus),
	.bondingout1(),
	.bondingout2(),
	.bondingout3(),
	.cfgaddlat(hmc_inst_CFGADDLAT_bus),
	.cfgbankaddrwidth(hmc_inst_CFGBANKADDRWIDTH_bus),
	.cfgcaswrlat(hmc_inst_CFGCASWRLAT_bus),
	.cfgcoladdrwidth(hmc_inst_CFGCOLADDRWIDTH_bus),
	.cfgcsaddrwidth(hmc_inst_CFGCSADDRWIDTH_bus),
	.cfgdevicewidth(hmc_inst_CFGDEVICEWIDTH_bus),
	.cfginterfacewidth(hmc_inst_CFGINTERFACEWIDTH_bus),
	.cfgrowaddrwidth(hmc_inst_CFGROWADDRWIDTH_bus),
	.cfgtcl(hmc_inst_CFGTCL_bus),
	.cfgtmrd(hmc_inst_CFGTMRD_bus),
	.cfgtrefi(hmc_inst_CFGTREFI_bus),
	.cfgtrfc(hmc_inst_CFGTRFC_bus),
	.cfgtwr(hmc_inst_CFGTWR_bus),
	.ctlcalbytelaneseln(),
	.ctlmemclkdisable(hmc_inst_CTLMEMCLKDISABLE_bus),
	.dramconfig(hmc_inst_DRAMCONFIG_bus),
	.mmrrdata(),
	.ordavstdata0(),
	.ordavstdata1(),
	.ordavstdata2(),
	.ordavstdata3(),
	.scrdata());
defparam hmc_inst.attr_counter_one_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_one_reset = "disabled";
defparam hmc_inst.attr_counter_zero_mask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_match = 64'b0000000000000000000000000000000000000000000000000000000000000000;
defparam hmc_inst.attr_counter_zero_reset = "disabled";
defparam hmc_inst.attr_debug_select_byte = 32'b00000000000000000000000000000000;
defparam hmc_inst.attr_static_config_valid = "disabled";
defparam hmc_inst.auto_pch_enable_0 = "disabled";
defparam hmc_inst.auto_pch_enable_1 = "disabled";
defparam hmc_inst.auto_pch_enable_2 = "disabled";
defparam hmc_inst.auto_pch_enable_3 = "disabled";
defparam hmc_inst.auto_pch_enable_4 = "disabled";
defparam hmc_inst.auto_pch_enable_5 = "disabled";
defparam hmc_inst.cal_req = "disabled";
defparam hmc_inst.cfg_burst_length = "bl_8";
defparam hmc_inst.cfg_interface_width = "dwidth_32";
defparam hmc_inst.cfg_self_rfsh_exit_cycles = "self_rfsh_exit_cycles_512";
defparam hmc_inst.cfg_starve_limit = "starve_limit_10";
defparam hmc_inst.cfg_type = "ddr3";
defparam hmc_inst.clr_intr = "no_clr_intr";
defparam hmc_inst.cmd_port_in_use_0 = "false";
defparam hmc_inst.cmd_port_in_use_1 = "false";
defparam hmc_inst.cmd_port_in_use_2 = "false";
defparam hmc_inst.cmd_port_in_use_3 = "false";
defparam hmc_inst.cmd_port_in_use_4 = "false";
defparam hmc_inst.cmd_port_in_use_5 = "false";
defparam hmc_inst.cport0_rdy_almost_full = "not_full";
defparam hmc_inst.cport0_rfifo_map = "fifo_0";
defparam hmc_inst.cport0_type = "disable";
defparam hmc_inst.cport0_wfifo_map = "fifo_0";
defparam hmc_inst.cport1_rdy_almost_full = "not_full";
defparam hmc_inst.cport1_rfifo_map = "fifo_0";
defparam hmc_inst.cport1_type = "disable";
defparam hmc_inst.cport1_wfifo_map = "fifo_0";
defparam hmc_inst.cport2_rdy_almost_full = "not_full";
defparam hmc_inst.cport2_rfifo_map = "fifo_0";
defparam hmc_inst.cport2_type = "disable";
defparam hmc_inst.cport2_wfifo_map = "fifo_0";
defparam hmc_inst.cport3_rdy_almost_full = "not_full";
defparam hmc_inst.cport3_rfifo_map = "fifo_0";
defparam hmc_inst.cport3_type = "disable";
defparam hmc_inst.cport3_wfifo_map = "fifo_0";
defparam hmc_inst.cport4_rdy_almost_full = "not_full";
defparam hmc_inst.cport4_rfifo_map = "fifo_0";
defparam hmc_inst.cport4_type = "disable";
defparam hmc_inst.cport4_wfifo_map = "fifo_0";
defparam hmc_inst.cport5_rdy_almost_full = "not_full";
defparam hmc_inst.cport5_rfifo_map = "fifo_0";
defparam hmc_inst.cport5_type = "disable";
defparam hmc_inst.cport5_wfifo_map = "fifo_0";
defparam hmc_inst.ctl_addr_order = "chip_row_bank_col";
defparam hmc_inst.ctl_ecc_enabled = "ctl_ecc_disabled";
defparam hmc_inst.ctl_ecc_rmw_enabled = "ctl_ecc_rmw_disabled";
defparam hmc_inst.ctl_regdimm_enabled = "regdimm_disabled";
defparam hmc_inst.ctl_usr_refresh = "ctl_usr_refresh_disabled";
defparam hmc_inst.ctrl_width = "data_width_64_bit";
defparam hmc_inst.cyc_to_rld_jars_0 = 1;
defparam hmc_inst.cyc_to_rld_jars_1 = 1;
defparam hmc_inst.cyc_to_rld_jars_2 = 1;
defparam hmc_inst.cyc_to_rld_jars_3 = 1;
defparam hmc_inst.cyc_to_rld_jars_4 = 1;
defparam hmc_inst.cyc_to_rld_jars_5 = 1;
defparam hmc_inst.delay_bonding = "bonding_latency_0";
defparam hmc_inst.dfx_bypass_enable = "dfx_bypass_disabled";
defparam hmc_inst.disable_merging = "merging_enabled";
defparam hmc_inst.ecc_dq_width = "ecc_dq_width_0";
defparam hmc_inst.enable_atpg = "disabled";
defparam hmc_inst.enable_bonding_0 = "disabled";
defparam hmc_inst.enable_bonding_1 = "disabled";
defparam hmc_inst.enable_bonding_2 = "disabled";
defparam hmc_inst.enable_bonding_3 = "disabled";
defparam hmc_inst.enable_bonding_4 = "disabled";
defparam hmc_inst.enable_bonding_5 = "disabled";
defparam hmc_inst.enable_bonding_wrapback = "disabled";
defparam hmc_inst.enable_burst_interrupt = "disabled";
defparam hmc_inst.enable_burst_terminate = "disabled";
defparam hmc_inst.enable_dqs_tracking = "enabled";
defparam hmc_inst.enable_ecc_code_overwrites = "disabled";
defparam hmc_inst.enable_fast_exit_ppd = "disabled";
defparam hmc_inst.enable_intr = "disabled";
defparam hmc_inst.enable_no_dm = "disabled";
defparam hmc_inst.enable_pipelineglobal = "disabled";
defparam hmc_inst.extra_ctl_clk_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_act_to_act_diff_bank = 0;
defparam hmc_inst.extra_ctl_clk_act_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_act_to_rdwr = 0;
defparam hmc_inst.extra_ctl_clk_arf_period = 0;
defparam hmc_inst.extra_ctl_clk_arf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_four_act_to_act = 0;
defparam hmc_inst.extra_ctl_clk_pch_all_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pch_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_pdn_period = 0;
defparam hmc_inst.extra_ctl_clk_pdn_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_rd_diff_chip = 0;
defparam hmc_inst.extra_ctl_clk_rd_to_wr = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_bc = 2;
defparam hmc_inst.extra_ctl_clk_rd_to_wr_diff_chip = 2;
defparam hmc_inst.extra_ctl_clk_srf_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_srf_to_zq_cal = 0;
defparam hmc_inst.extra_ctl_clk_wr_ap_to_valid = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_pch = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_rd = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_bc = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_rd_diff_chip = 3;
defparam hmc_inst.extra_ctl_clk_wr_to_wr = 0;
defparam hmc_inst.extra_ctl_clk_wr_to_wr_diff_chip = 0;
defparam hmc_inst.gen_dbe = "gen_dbe_disabled";
defparam hmc_inst.gen_sbe = "gen_sbe_disabled";
defparam hmc_inst.inc_sync = "fifo_set_2";
defparam hmc_inst.local_if_cs_width = "addr_width_0";
defparam hmc_inst.mask_corr_dropped_intr = "disabled";
defparam hmc_inst.mask_dbe_intr = "disabled";
defparam hmc_inst.mask_sbe_intr = "disabled";
defparam hmc_inst.mem_auto_pd_cycles = 0;
defparam hmc_inst.mem_clk_entry_cycles = 10;
defparam hmc_inst.mem_if_al = "al_0";
defparam hmc_inst.mem_if_bankaddr_width = "addr_width_3";
defparam hmc_inst.mem_if_burstlength = "mem_if_burstlength_8";
defparam hmc_inst.mem_if_coladdr_width = "addr_width_10";
defparam hmc_inst.mem_if_cs_per_rank = "mem_if_cs_per_rank_1";
defparam hmc_inst.mem_if_cs_width = "mem_if_cs_width_1";
defparam hmc_inst.mem_if_dq_per_chip = "mem_if_dq_per_chip_8";
defparam hmc_inst.mem_if_dqs_width = "dqs_width_4";
defparam hmc_inst.mem_if_dwidth = "mem_if_dwidth_32";
defparam hmc_inst.mem_if_memtype = "ddr3_sdram";
defparam hmc_inst.mem_if_rowaddr_width = "addr_width_15";
defparam hmc_inst.mem_if_speedbin = "ddr3_1600_8_8_8";
defparam hmc_inst.mem_if_tccd = "tccd_4";
defparam hmc_inst.mem_if_tcl = "tcl_7";
defparam hmc_inst.mem_if_tcwl = "tcwl_7";
defparam hmc_inst.mem_if_tfaw = "tfaw_18";
defparam hmc_inst.mem_if_tmrd = "tmrd_4";
defparam hmc_inst.mem_if_tras = "tras_15";
defparam hmc_inst.mem_if_trc = "trc_20";
defparam hmc_inst.mem_if_trcd = "trcd_6";
defparam hmc_inst.mem_if_trefi = 3120;
defparam hmc_inst.mem_if_trfc = 120;
defparam hmc_inst.mem_if_trp = "trp_6";
defparam hmc_inst.mem_if_trrd = "trrd_3";
defparam hmc_inst.mem_if_trtp = "trtp_3";
defparam hmc_inst.mem_if_twr = "twr_6";
defparam hmc_inst.mem_if_twtr = "twtr_4";
defparam hmc_inst.mmr_cfg_mem_bl = "mp_bl_8";
defparam hmc_inst.output_regd = "disabled";
defparam hmc_inst.pdn_exit_cycles = "slow_exit";
defparam hmc_inst.port0_width = "port_32_bit";
defparam hmc_inst.port1_width = "port_32_bit";
defparam hmc_inst.port2_width = "port_32_bit";
defparam hmc_inst.port3_width = "port_32_bit";
defparam hmc_inst.port4_width = "port_32_bit";
defparam hmc_inst.port5_width = "port_32_bit";
defparam hmc_inst.power_saving_exit_cycles = 5;
defparam hmc_inst.priority_0_0 = "weight_0";
defparam hmc_inst.priority_0_1 = "weight_0";
defparam hmc_inst.priority_0_2 = "weight_0";
defparam hmc_inst.priority_0_3 = "weight_0";
defparam hmc_inst.priority_0_4 = "weight_0";
defparam hmc_inst.priority_0_5 = "weight_0";
defparam hmc_inst.priority_1_0 = "weight_0";
defparam hmc_inst.priority_1_1 = "weight_0";
defparam hmc_inst.priority_1_2 = "weight_0";
defparam hmc_inst.priority_1_3 = "weight_0";
defparam hmc_inst.priority_1_4 = "weight_0";
defparam hmc_inst.priority_1_5 = "weight_0";
defparam hmc_inst.priority_2_0 = "weight_0";
defparam hmc_inst.priority_2_1 = "weight_0";
defparam hmc_inst.priority_2_2 = "weight_0";
defparam hmc_inst.priority_2_3 = "weight_0";
defparam hmc_inst.priority_2_4 = "weight_0";
defparam hmc_inst.priority_2_5 = "weight_0";
defparam hmc_inst.priority_3_0 = "weight_0";
defparam hmc_inst.priority_3_1 = "weight_0";
defparam hmc_inst.priority_3_2 = "weight_0";
defparam hmc_inst.priority_3_3 = "weight_0";
defparam hmc_inst.priority_3_4 = "weight_0";
defparam hmc_inst.priority_3_5 = "weight_0";
defparam hmc_inst.priority_4_0 = "weight_0";
defparam hmc_inst.priority_4_1 = "weight_0";
defparam hmc_inst.priority_4_2 = "weight_0";
defparam hmc_inst.priority_4_3 = "weight_0";
defparam hmc_inst.priority_4_4 = "weight_0";
defparam hmc_inst.priority_4_5 = "weight_0";
defparam hmc_inst.priority_5_0 = "weight_0";
defparam hmc_inst.priority_5_1 = "weight_0";
defparam hmc_inst.priority_5_2 = "weight_0";
defparam hmc_inst.priority_5_3 = "weight_0";
defparam hmc_inst.priority_5_4 = "weight_0";
defparam hmc_inst.priority_5_5 = "weight_0";
defparam hmc_inst.priority_6_0 = "weight_0";
defparam hmc_inst.priority_6_1 = "weight_0";
defparam hmc_inst.priority_6_2 = "weight_0";
defparam hmc_inst.priority_6_3 = "weight_0";
defparam hmc_inst.priority_6_4 = "weight_0";
defparam hmc_inst.priority_6_5 = "weight_0";
defparam hmc_inst.priority_7_0 = "weight_0";
defparam hmc_inst.priority_7_1 = "weight_0";
defparam hmc_inst.priority_7_2 = "weight_0";
defparam hmc_inst.priority_7_3 = "weight_0";
defparam hmc_inst.priority_7_4 = "weight_0";
defparam hmc_inst.priority_7_5 = "weight_0";
defparam hmc_inst.priority_remap = 0;
defparam hmc_inst.rcfg_static_weight_0 = "weight_0";
defparam hmc_inst.rcfg_static_weight_1 = "weight_0";
defparam hmc_inst.rcfg_static_weight_2 = "weight_0";
defparam hmc_inst.rcfg_static_weight_3 = "weight_0";
defparam hmc_inst.rcfg_static_weight_4 = "weight_0";
defparam hmc_inst.rcfg_static_weight_5 = "weight_0";
defparam hmc_inst.rcfg_sum_wt_priority_0 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_1 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_2 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_3 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_4 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_5 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_6 = 0;
defparam hmc_inst.rcfg_sum_wt_priority_7 = 0;
defparam hmc_inst.rcfg_user_priority_0 = "priority_1";
defparam hmc_inst.rcfg_user_priority_1 = "priority_1";
defparam hmc_inst.rcfg_user_priority_2 = "priority_1";
defparam hmc_inst.rcfg_user_priority_3 = "priority_1";
defparam hmc_inst.rcfg_user_priority_4 = "priority_1";
defparam hmc_inst.rcfg_user_priority_5 = "priority_1";
defparam hmc_inst.rd_dwidth_0 = "dwidth_0";
defparam hmc_inst.rd_dwidth_1 = "dwidth_0";
defparam hmc_inst.rd_dwidth_2 = "dwidth_0";
defparam hmc_inst.rd_dwidth_3 = "dwidth_0";
defparam hmc_inst.rd_dwidth_4 = "dwidth_0";
defparam hmc_inst.rd_dwidth_5 = "dwidth_0";
defparam hmc_inst.rd_fifo_in_use_0 = "false";
defparam hmc_inst.rd_fifo_in_use_1 = "false";
defparam hmc_inst.rd_fifo_in_use_2 = "false";
defparam hmc_inst.rd_fifo_in_use_3 = "false";
defparam hmc_inst.rd_port_info_0 = "use_no";
defparam hmc_inst.rd_port_info_1 = "use_no";
defparam hmc_inst.rd_port_info_2 = "use_no";
defparam hmc_inst.rd_port_info_3 = "use_no";
defparam hmc_inst.rd_port_info_4 = "use_no";
defparam hmc_inst.rd_port_info_5 = "use_no";
defparam hmc_inst.read_odt_chip = "odt_disabled";
defparam hmc_inst.reorder_data = "data_reordering";
defparam hmc_inst.rfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.rfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.single_ready_0 = "concatenate_rdy";
defparam hmc_inst.single_ready_1 = "concatenate_rdy";
defparam hmc_inst.single_ready_2 = "concatenate_rdy";
defparam hmc_inst.single_ready_3 = "concatenate_rdy";
defparam hmc_inst.static_weight_0 = "weight_0";
defparam hmc_inst.static_weight_1 = "weight_0";
defparam hmc_inst.static_weight_2 = "weight_0";
defparam hmc_inst.static_weight_3 = "weight_0";
defparam hmc_inst.static_weight_4 = "weight_0";
defparam hmc_inst.static_weight_5 = "weight_0";
defparam hmc_inst.sum_wt_priority_0 = 0;
defparam hmc_inst.sum_wt_priority_1 = 0;
defparam hmc_inst.sum_wt_priority_2 = 0;
defparam hmc_inst.sum_wt_priority_3 = 0;
defparam hmc_inst.sum_wt_priority_4 = 0;
defparam hmc_inst.sum_wt_priority_5 = 0;
defparam hmc_inst.sum_wt_priority_6 = 0;
defparam hmc_inst.sum_wt_priority_7 = 0;
defparam hmc_inst.sync_mode_0 = "asynchronous";
defparam hmc_inst.sync_mode_1 = "asynchronous";
defparam hmc_inst.sync_mode_2 = "asynchronous";
defparam hmc_inst.sync_mode_3 = "asynchronous";
defparam hmc_inst.sync_mode_4 = "asynchronous";
defparam hmc_inst.sync_mode_5 = "asynchronous";
defparam hmc_inst.test_mode = "normal_mode";
defparam hmc_inst.thld_jar1_0 = "threshold_32";
defparam hmc_inst.thld_jar1_1 = "threshold_32";
defparam hmc_inst.thld_jar1_2 = "threshold_32";
defparam hmc_inst.thld_jar1_3 = "threshold_32";
defparam hmc_inst.thld_jar1_4 = "threshold_32";
defparam hmc_inst.thld_jar1_5 = "threshold_32";
defparam hmc_inst.thld_jar2_0 = "threshold_16";
defparam hmc_inst.thld_jar2_1 = "threshold_16";
defparam hmc_inst.thld_jar2_2 = "threshold_16";
defparam hmc_inst.thld_jar2_3 = "threshold_16";
defparam hmc_inst.thld_jar2_4 = "threshold_16";
defparam hmc_inst.thld_jar2_5 = "threshold_16";
defparam hmc_inst.use_almost_empty_0 = "empty";
defparam hmc_inst.use_almost_empty_1 = "empty";
defparam hmc_inst.use_almost_empty_2 = "empty";
defparam hmc_inst.use_almost_empty_3 = "empty";
defparam hmc_inst.user_ecc_en = "disable";
defparam hmc_inst.user_priority_0 = "priority_1";
defparam hmc_inst.user_priority_1 = "priority_1";
defparam hmc_inst.user_priority_2 = "priority_1";
defparam hmc_inst.user_priority_3 = "priority_1";
defparam hmc_inst.user_priority_4 = "priority_1";
defparam hmc_inst.user_priority_5 = "priority_1";
defparam hmc_inst.wfifo0_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo0_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo1_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo1_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo2_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo2_rdy_almost_full = "not_full";
defparam hmc_inst.wfifo3_cport_map = "cmd_port_0";
defparam hmc_inst.wfifo3_rdy_almost_full = "not_full";
defparam hmc_inst.wr_dwidth_0 = "dwidth_0";
defparam hmc_inst.wr_dwidth_1 = "dwidth_0";
defparam hmc_inst.wr_dwidth_2 = "dwidth_0";
defparam hmc_inst.wr_dwidth_3 = "dwidth_0";
defparam hmc_inst.wr_dwidth_4 = "dwidth_0";
defparam hmc_inst.wr_dwidth_5 = "dwidth_0";
defparam hmc_inst.wr_fifo_in_use_0 = "false";
defparam hmc_inst.wr_fifo_in_use_1 = "false";
defparam hmc_inst.wr_fifo_in_use_2 = "false";
defparam hmc_inst.wr_fifo_in_use_3 = "false";
defparam hmc_inst.wr_port_info_0 = "use_no";
defparam hmc_inst.wr_port_info_1 = "use_no";
defparam hmc_inst.wr_port_info_2 = "use_no";
defparam hmc_inst.wr_port_info_3 = "use_no";
defparam hmc_inst.wr_port_info_4 = "use_no";
defparam hmc_inst.wr_port_info_5 = "use_no";
defparam hmc_inst.write_odt_chip = "write_chip0_odt0_chip1";

endmodule

module terminal_qsys_altera_mem_if_oct_cyclonev (
	parallelterminationcontrol,
	seriesterminationcontrol,
	oct_rzqin)/* synthesis synthesis_greybox=0 */;
output 	[15:0] parallelterminationcontrol;
output 	[15:0] seriesterminationcontrol;
input 	oct_rzqin;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sd1a_0~O_CLKUSRDFTOUT ;
wire \wire_sd1a_serdataout[0] ;

wire [15:0] sd2a_0_PARALLELTERMINATIONCONTROL_bus;
wire [15:0] sd2a_0_SERIESTERMINATIONCONTROL_bus;

assign parallelterminationcontrol[0] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[0];
assign parallelterminationcontrol[1] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[1];
assign parallelterminationcontrol[2] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[2];
assign parallelterminationcontrol[3] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[3];
assign parallelterminationcontrol[4] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[4];
assign parallelterminationcontrol[5] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[5];
assign parallelterminationcontrol[6] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[6];
assign parallelterminationcontrol[7] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[7];
assign parallelterminationcontrol[8] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[8];
assign parallelterminationcontrol[9] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[9];
assign parallelterminationcontrol[10] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[10];
assign parallelterminationcontrol[11] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[11];
assign parallelterminationcontrol[12] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[12];
assign parallelterminationcontrol[13] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[13];
assign parallelterminationcontrol[14] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[14];
assign parallelterminationcontrol[15] = sd2a_0_PARALLELTERMINATIONCONTROL_bus[15];

assign seriesterminationcontrol[0] = sd2a_0_SERIESTERMINATIONCONTROL_bus[0];
assign seriesterminationcontrol[1] = sd2a_0_SERIESTERMINATIONCONTROL_bus[1];
assign seriesterminationcontrol[2] = sd2a_0_SERIESTERMINATIONCONTROL_bus[2];
assign seriesterminationcontrol[3] = sd2a_0_SERIESTERMINATIONCONTROL_bus[3];
assign seriesterminationcontrol[4] = sd2a_0_SERIESTERMINATIONCONTROL_bus[4];
assign seriesterminationcontrol[5] = sd2a_0_SERIESTERMINATIONCONTROL_bus[5];
assign seriesterminationcontrol[6] = sd2a_0_SERIESTERMINATIONCONTROL_bus[6];
assign seriesterminationcontrol[7] = sd2a_0_SERIESTERMINATIONCONTROL_bus[7];
assign seriesterminationcontrol[8] = sd2a_0_SERIESTERMINATIONCONTROL_bus[8];
assign seriesterminationcontrol[9] = sd2a_0_SERIESTERMINATIONCONTROL_bus[9];
assign seriesterminationcontrol[10] = sd2a_0_SERIESTERMINATIONCONTROL_bus[10];
assign seriesterminationcontrol[11] = sd2a_0_SERIESTERMINATIONCONTROL_bus[11];
assign seriesterminationcontrol[12] = sd2a_0_SERIESTERMINATIONCONTROL_bus[12];
assign seriesterminationcontrol[13] = sd2a_0_SERIESTERMINATIONCONTROL_bus[13];
assign seriesterminationcontrol[14] = sd2a_0_SERIESTERMINATIONCONTROL_bus[14];
assign seriesterminationcontrol[15] = sd2a_0_SERIESTERMINATIONCONTROL_bus[15];

cyclonev_termination_logic sd2a_0(
	.s2pload(gnd),
	.scanclk(gnd),
	.scanenable(gnd),
	.serdata(\wire_sd1a_serdataout[0] ),
	.enser(4'b0000),
	.parallelterminationcontrol(sd2a_0_PARALLELTERMINATIONCONTROL_bus),
	.seriesterminationcontrol(sd2a_0_SERIESTERMINATIONCONTROL_bus));

cyclonev_termination sd1a_0(
	.clkenusr(gnd),
	.clkusr(gnd),
	.enserusr(gnd),
	.nclrusr(gnd),
	.rzqin(oct_rzqin),
	.scanclk(gnd),
	.scanen(gnd),
	.scanin(gnd),
	.serdatafromcore(gnd),
	.serdatain(gnd),
	.otherenser(10'b0000000000),
	.clkusrdftout(\sd1a_0~O_CLKUSRDFTOUT ),
	.compoutrdn(),
	.compoutrup(),
	.enserout(),
	.scanout(),
	.serdataout(\wire_sd1a_serdataout[0] ),
	.serdatatocore());

endmodule

module terminal_qsys_hps_sdram_p0 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid_0,
	ctl_reset_n,
	afi_rdata_0,
	afi_rdata_1,
	afi_rdata_2,
	afi_rdata_3,
	afi_rdata_4,
	afi_rdata_5,
	afi_rdata_6,
	afi_rdata_7,
	afi_rdata_8,
	afi_rdata_9,
	afi_rdata_10,
	afi_rdata_11,
	afi_rdata_12,
	afi_rdata_13,
	afi_rdata_14,
	afi_rdata_15,
	afi_rdata_16,
	afi_rdata_17,
	afi_rdata_18,
	afi_rdata_19,
	afi_rdata_20,
	afi_rdata_21,
	afi_rdata_22,
	afi_rdata_23,
	afi_rdata_24,
	afi_rdata_25,
	afi_rdata_26,
	afi_rdata_27,
	afi_rdata_28,
	afi_rdata_29,
	afi_rdata_30,
	afi_rdata_31,
	afi_rdata_32,
	afi_rdata_33,
	afi_rdata_34,
	afi_rdata_35,
	afi_rdata_36,
	afi_rdata_37,
	afi_rdata_38,
	afi_rdata_39,
	afi_rdata_40,
	afi_rdata_41,
	afi_rdata_42,
	afi_rdata_43,
	afi_rdata_44,
	afi_rdata_45,
	afi_rdata_46,
	afi_rdata_47,
	afi_rdata_48,
	afi_rdata_49,
	afi_rdata_50,
	afi_rdata_51,
	afi_rdata_52,
	afi_rdata_53,
	afi_rdata_54,
	afi_rdata_55,
	afi_rdata_56,
	afi_rdata_57,
	afi_rdata_58,
	afi_rdata_59,
	afi_rdata_60,
	afi_rdata_61,
	afi_rdata_62,
	afi_rdata_63,
	afi_rdata_64,
	afi_rdata_65,
	afi_rdata_66,
	afi_rdata_67,
	afi_rdata_68,
	afi_rdata_69,
	afi_rdata_70,
	afi_rdata_71,
	afi_rdata_72,
	afi_rdata_73,
	afi_rdata_74,
	afi_rdata_75,
	afi_rdata_76,
	afi_rdata_77,
	afi_rdata_78,
	afi_rdata_79,
	afi_wlat_0,
	afi_wlat_1,
	afi_wlat_2,
	afi_wlat_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n_0,
	afi_ras_n_0,
	afi_rst_n_0,
	afi_we_n_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_addr_14,
	afi_addr_15,
	afi_addr_16,
	afi_addr_17,
	afi_addr_18,
	afi_addr_19,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_cke_0,
	afi_cke_1,
	afi_cs_n_0,
	afi_cs_n_1,
	afi_dm_int_0,
	afi_dm_int_1,
	afi_dm_int_2,
	afi_dm_int_3,
	afi_dm_int_4,
	afi_dm_int_5,
	afi_dm_int_6,
	afi_dm_int_7,
	afi_dm_int_8,
	afi_dm_int_9,
	afi_dqs_burst_0,
	afi_dqs_burst_1,
	afi_dqs_burst_2,
	afi_dqs_burst_3,
	afi_dqs_burst_4,
	afi_odt_0,
	afi_odt_1,
	afi_rdata_en_0,
	afi_rdata_en_1,
	afi_rdata_en_2,
	afi_rdata_en_3,
	afi_rdata_en_4,
	afi_rdata_en_full_0,
	afi_rdata_en_full_1,
	afi_rdata_en_full_2,
	afi_rdata_en_full_3,
	afi_rdata_en_full_4,
	afi_wdata_int_0,
	afi_wdata_int_1,
	afi_wdata_int_2,
	afi_wdata_int_3,
	afi_wdata_int_4,
	afi_wdata_int_5,
	afi_wdata_int_6,
	afi_wdata_int_7,
	afi_wdata_int_8,
	afi_wdata_int_9,
	afi_wdata_int_10,
	afi_wdata_int_11,
	afi_wdata_int_12,
	afi_wdata_int_13,
	afi_wdata_int_14,
	afi_wdata_int_15,
	afi_wdata_int_16,
	afi_wdata_int_17,
	afi_wdata_int_18,
	afi_wdata_int_19,
	afi_wdata_int_20,
	afi_wdata_int_21,
	afi_wdata_int_22,
	afi_wdata_int_23,
	afi_wdata_int_24,
	afi_wdata_int_25,
	afi_wdata_int_26,
	afi_wdata_int_27,
	afi_wdata_int_28,
	afi_wdata_int_29,
	afi_wdata_int_30,
	afi_wdata_int_31,
	afi_wdata_int_32,
	afi_wdata_int_33,
	afi_wdata_int_34,
	afi_wdata_int_35,
	afi_wdata_int_36,
	afi_wdata_int_37,
	afi_wdata_int_38,
	afi_wdata_int_39,
	afi_wdata_int_40,
	afi_wdata_int_41,
	afi_wdata_int_42,
	afi_wdata_int_43,
	afi_wdata_int_44,
	afi_wdata_int_45,
	afi_wdata_int_46,
	afi_wdata_int_47,
	afi_wdata_int_48,
	afi_wdata_int_49,
	afi_wdata_int_50,
	afi_wdata_int_51,
	afi_wdata_int_52,
	afi_wdata_int_53,
	afi_wdata_int_54,
	afi_wdata_int_55,
	afi_wdata_int_56,
	afi_wdata_int_57,
	afi_wdata_int_58,
	afi_wdata_int_59,
	afi_wdata_int_60,
	afi_wdata_int_61,
	afi_wdata_int_62,
	afi_wdata_int_63,
	afi_wdata_int_64,
	afi_wdata_int_65,
	afi_wdata_int_66,
	afi_wdata_int_67,
	afi_wdata_int_68,
	afi_wdata_int_69,
	afi_wdata_int_70,
	afi_wdata_int_71,
	afi_wdata_int_72,
	afi_wdata_int_73,
	afi_wdata_int_74,
	afi_wdata_int_75,
	afi_wdata_int_76,
	afi_wdata_int_77,
	afi_wdata_int_78,
	afi_wdata_int_79,
	afi_wdata_valid_0,
	afi_wdata_valid_1,
	afi_wdata_valid_2,
	afi_wdata_valid_3,
	afi_wdata_valid_4,
	cfg_addlat_wire_0,
	cfg_addlat_wire_1,
	cfg_addlat_wire_2,
	cfg_addlat_wire_3,
	cfg_addlat_wire_4,
	cfg_bankaddrwidth_wire_0,
	cfg_bankaddrwidth_wire_1,
	cfg_bankaddrwidth_wire_2,
	cfg_caswrlat_wire_0,
	cfg_caswrlat_wire_1,
	cfg_caswrlat_wire_2,
	cfg_caswrlat_wire_3,
	cfg_coladdrwidth_wire_0,
	cfg_coladdrwidth_wire_1,
	cfg_coladdrwidth_wire_2,
	cfg_coladdrwidth_wire_3,
	cfg_coladdrwidth_wire_4,
	cfg_csaddrwidth_wire_0,
	cfg_csaddrwidth_wire_1,
	cfg_csaddrwidth_wire_2,
	cfg_devicewidth_wire_0,
	cfg_devicewidth_wire_1,
	cfg_devicewidth_wire_2,
	cfg_devicewidth_wire_3,
	cfg_interfacewidth_wire_0,
	cfg_interfacewidth_wire_1,
	cfg_interfacewidth_wire_2,
	cfg_interfacewidth_wire_3,
	cfg_interfacewidth_wire_4,
	cfg_interfacewidth_wire_5,
	cfg_interfacewidth_wire_6,
	cfg_interfacewidth_wire_7,
	cfg_rowaddrwidth_wire_0,
	cfg_rowaddrwidth_wire_1,
	cfg_rowaddrwidth_wire_2,
	cfg_rowaddrwidth_wire_3,
	cfg_rowaddrwidth_wire_4,
	cfg_tcl_wire_0,
	cfg_tcl_wire_1,
	cfg_tcl_wire_2,
	cfg_tcl_wire_3,
	cfg_tcl_wire_4,
	cfg_tmrd_wire_0,
	cfg_tmrd_wire_1,
	cfg_tmrd_wire_2,
	cfg_tmrd_wire_3,
	cfg_trefi_wire_0,
	cfg_trefi_wire_1,
	cfg_trefi_wire_2,
	cfg_trefi_wire_3,
	cfg_trefi_wire_4,
	cfg_trefi_wire_5,
	cfg_trefi_wire_6,
	cfg_trefi_wire_7,
	cfg_trefi_wire_8,
	cfg_trefi_wire_9,
	cfg_trefi_wire_10,
	cfg_trefi_wire_11,
	cfg_trefi_wire_12,
	cfg_trfc_wire_0,
	cfg_trfc_wire_1,
	cfg_trfc_wire_2,
	cfg_trfc_wire_3,
	cfg_trfc_wire_4,
	cfg_trfc_wire_5,
	cfg_trfc_wire_6,
	cfg_trfc_wire_7,
	cfg_twr_wire_0,
	cfg_twr_wire_1,
	cfg_twr_wire_2,
	cfg_twr_wire_3,
	afi_mem_clk_disable_0,
	cfg_dramconfig_wire_0,
	cfg_dramconfig_wire_1,
	cfg_dramconfig_wire_2,
	cfg_dramconfig_wire_3,
	cfg_dramconfig_wire_4,
	cfg_dramconfig_wire_5,
	cfg_dramconfig_wire_6,
	cfg_dramconfig_wire_7,
	cfg_dramconfig_wire_8,
	cfg_dramconfig_wire_9,
	cfg_dramconfig_wire_10,
	cfg_dramconfig_wire_11,
	cfg_dramconfig_wire_12,
	cfg_dramconfig_wire_13,
	cfg_dramconfig_wire_14,
	cfg_dramconfig_wire_15,
	cfg_dramconfig_wire_16,
	cfg_dramconfig_wire_17,
	cfg_dramconfig_wire_18,
	cfg_dramconfig_wire_19,
	cfg_dramconfig_wire_20,
	ctl_clk,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	afi_rdata_valid_0;
output 	ctl_reset_n;
output 	afi_rdata_0;
output 	afi_rdata_1;
output 	afi_rdata_2;
output 	afi_rdata_3;
output 	afi_rdata_4;
output 	afi_rdata_5;
output 	afi_rdata_6;
output 	afi_rdata_7;
output 	afi_rdata_8;
output 	afi_rdata_9;
output 	afi_rdata_10;
output 	afi_rdata_11;
output 	afi_rdata_12;
output 	afi_rdata_13;
output 	afi_rdata_14;
output 	afi_rdata_15;
output 	afi_rdata_16;
output 	afi_rdata_17;
output 	afi_rdata_18;
output 	afi_rdata_19;
output 	afi_rdata_20;
output 	afi_rdata_21;
output 	afi_rdata_22;
output 	afi_rdata_23;
output 	afi_rdata_24;
output 	afi_rdata_25;
output 	afi_rdata_26;
output 	afi_rdata_27;
output 	afi_rdata_28;
output 	afi_rdata_29;
output 	afi_rdata_30;
output 	afi_rdata_31;
output 	afi_rdata_32;
output 	afi_rdata_33;
output 	afi_rdata_34;
output 	afi_rdata_35;
output 	afi_rdata_36;
output 	afi_rdata_37;
output 	afi_rdata_38;
output 	afi_rdata_39;
output 	afi_rdata_40;
output 	afi_rdata_41;
output 	afi_rdata_42;
output 	afi_rdata_43;
output 	afi_rdata_44;
output 	afi_rdata_45;
output 	afi_rdata_46;
output 	afi_rdata_47;
output 	afi_rdata_48;
output 	afi_rdata_49;
output 	afi_rdata_50;
output 	afi_rdata_51;
output 	afi_rdata_52;
output 	afi_rdata_53;
output 	afi_rdata_54;
output 	afi_rdata_55;
output 	afi_rdata_56;
output 	afi_rdata_57;
output 	afi_rdata_58;
output 	afi_rdata_59;
output 	afi_rdata_60;
output 	afi_rdata_61;
output 	afi_rdata_62;
output 	afi_rdata_63;
output 	afi_rdata_64;
output 	afi_rdata_65;
output 	afi_rdata_66;
output 	afi_rdata_67;
output 	afi_rdata_68;
output 	afi_rdata_69;
output 	afi_rdata_70;
output 	afi_rdata_71;
output 	afi_rdata_72;
output 	afi_rdata_73;
output 	afi_rdata_74;
output 	afi_rdata_75;
output 	afi_rdata_76;
output 	afi_rdata_77;
output 	afi_rdata_78;
output 	afi_rdata_79;
output 	afi_wlat_0;
output 	afi_wlat_1;
output 	afi_wlat_2;
output 	afi_wlat_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	afi_cas_n_0;
input 	afi_ras_n_0;
input 	afi_rst_n_0;
input 	afi_we_n_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_addr_14;
input 	afi_addr_15;
input 	afi_addr_16;
input 	afi_addr_17;
input 	afi_addr_18;
input 	afi_addr_19;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_cke_0;
input 	afi_cke_1;
input 	afi_cs_n_0;
input 	afi_cs_n_1;
input 	afi_dm_int_0;
input 	afi_dm_int_1;
input 	afi_dm_int_2;
input 	afi_dm_int_3;
input 	afi_dm_int_4;
input 	afi_dm_int_5;
input 	afi_dm_int_6;
input 	afi_dm_int_7;
input 	afi_dm_int_8;
input 	afi_dm_int_9;
input 	afi_dqs_burst_0;
input 	afi_dqs_burst_1;
input 	afi_dqs_burst_2;
input 	afi_dqs_burst_3;
input 	afi_dqs_burst_4;
input 	afi_odt_0;
input 	afi_odt_1;
input 	afi_rdata_en_0;
input 	afi_rdata_en_1;
input 	afi_rdata_en_2;
input 	afi_rdata_en_3;
input 	afi_rdata_en_4;
input 	afi_rdata_en_full_0;
input 	afi_rdata_en_full_1;
input 	afi_rdata_en_full_2;
input 	afi_rdata_en_full_3;
input 	afi_rdata_en_full_4;
input 	afi_wdata_int_0;
input 	afi_wdata_int_1;
input 	afi_wdata_int_2;
input 	afi_wdata_int_3;
input 	afi_wdata_int_4;
input 	afi_wdata_int_5;
input 	afi_wdata_int_6;
input 	afi_wdata_int_7;
input 	afi_wdata_int_8;
input 	afi_wdata_int_9;
input 	afi_wdata_int_10;
input 	afi_wdata_int_11;
input 	afi_wdata_int_12;
input 	afi_wdata_int_13;
input 	afi_wdata_int_14;
input 	afi_wdata_int_15;
input 	afi_wdata_int_16;
input 	afi_wdata_int_17;
input 	afi_wdata_int_18;
input 	afi_wdata_int_19;
input 	afi_wdata_int_20;
input 	afi_wdata_int_21;
input 	afi_wdata_int_22;
input 	afi_wdata_int_23;
input 	afi_wdata_int_24;
input 	afi_wdata_int_25;
input 	afi_wdata_int_26;
input 	afi_wdata_int_27;
input 	afi_wdata_int_28;
input 	afi_wdata_int_29;
input 	afi_wdata_int_30;
input 	afi_wdata_int_31;
input 	afi_wdata_int_32;
input 	afi_wdata_int_33;
input 	afi_wdata_int_34;
input 	afi_wdata_int_35;
input 	afi_wdata_int_36;
input 	afi_wdata_int_37;
input 	afi_wdata_int_38;
input 	afi_wdata_int_39;
input 	afi_wdata_int_40;
input 	afi_wdata_int_41;
input 	afi_wdata_int_42;
input 	afi_wdata_int_43;
input 	afi_wdata_int_44;
input 	afi_wdata_int_45;
input 	afi_wdata_int_46;
input 	afi_wdata_int_47;
input 	afi_wdata_int_48;
input 	afi_wdata_int_49;
input 	afi_wdata_int_50;
input 	afi_wdata_int_51;
input 	afi_wdata_int_52;
input 	afi_wdata_int_53;
input 	afi_wdata_int_54;
input 	afi_wdata_int_55;
input 	afi_wdata_int_56;
input 	afi_wdata_int_57;
input 	afi_wdata_int_58;
input 	afi_wdata_int_59;
input 	afi_wdata_int_60;
input 	afi_wdata_int_61;
input 	afi_wdata_int_62;
input 	afi_wdata_int_63;
input 	afi_wdata_int_64;
input 	afi_wdata_int_65;
input 	afi_wdata_int_66;
input 	afi_wdata_int_67;
input 	afi_wdata_int_68;
input 	afi_wdata_int_69;
input 	afi_wdata_int_70;
input 	afi_wdata_int_71;
input 	afi_wdata_int_72;
input 	afi_wdata_int_73;
input 	afi_wdata_int_74;
input 	afi_wdata_int_75;
input 	afi_wdata_int_76;
input 	afi_wdata_int_77;
input 	afi_wdata_int_78;
input 	afi_wdata_int_79;
input 	afi_wdata_valid_0;
input 	afi_wdata_valid_1;
input 	afi_wdata_valid_2;
input 	afi_wdata_valid_3;
input 	afi_wdata_valid_4;
input 	cfg_addlat_wire_0;
input 	cfg_addlat_wire_1;
input 	cfg_addlat_wire_2;
input 	cfg_addlat_wire_3;
input 	cfg_addlat_wire_4;
input 	cfg_bankaddrwidth_wire_0;
input 	cfg_bankaddrwidth_wire_1;
input 	cfg_bankaddrwidth_wire_2;
input 	cfg_caswrlat_wire_0;
input 	cfg_caswrlat_wire_1;
input 	cfg_caswrlat_wire_2;
input 	cfg_caswrlat_wire_3;
input 	cfg_coladdrwidth_wire_0;
input 	cfg_coladdrwidth_wire_1;
input 	cfg_coladdrwidth_wire_2;
input 	cfg_coladdrwidth_wire_3;
input 	cfg_coladdrwidth_wire_4;
input 	cfg_csaddrwidth_wire_0;
input 	cfg_csaddrwidth_wire_1;
input 	cfg_csaddrwidth_wire_2;
input 	cfg_devicewidth_wire_0;
input 	cfg_devicewidth_wire_1;
input 	cfg_devicewidth_wire_2;
input 	cfg_devicewidth_wire_3;
input 	cfg_interfacewidth_wire_0;
input 	cfg_interfacewidth_wire_1;
input 	cfg_interfacewidth_wire_2;
input 	cfg_interfacewidth_wire_3;
input 	cfg_interfacewidth_wire_4;
input 	cfg_interfacewidth_wire_5;
input 	cfg_interfacewidth_wire_6;
input 	cfg_interfacewidth_wire_7;
input 	cfg_rowaddrwidth_wire_0;
input 	cfg_rowaddrwidth_wire_1;
input 	cfg_rowaddrwidth_wire_2;
input 	cfg_rowaddrwidth_wire_3;
input 	cfg_rowaddrwidth_wire_4;
input 	cfg_tcl_wire_0;
input 	cfg_tcl_wire_1;
input 	cfg_tcl_wire_2;
input 	cfg_tcl_wire_3;
input 	cfg_tcl_wire_4;
input 	cfg_tmrd_wire_0;
input 	cfg_tmrd_wire_1;
input 	cfg_tmrd_wire_2;
input 	cfg_tmrd_wire_3;
input 	cfg_trefi_wire_0;
input 	cfg_trefi_wire_1;
input 	cfg_trefi_wire_2;
input 	cfg_trefi_wire_3;
input 	cfg_trefi_wire_4;
input 	cfg_trefi_wire_5;
input 	cfg_trefi_wire_6;
input 	cfg_trefi_wire_7;
input 	cfg_trefi_wire_8;
input 	cfg_trefi_wire_9;
input 	cfg_trefi_wire_10;
input 	cfg_trefi_wire_11;
input 	cfg_trefi_wire_12;
input 	cfg_trfc_wire_0;
input 	cfg_trfc_wire_1;
input 	cfg_trfc_wire_2;
input 	cfg_trfc_wire_3;
input 	cfg_trfc_wire_4;
input 	cfg_trfc_wire_5;
input 	cfg_trfc_wire_6;
input 	cfg_trfc_wire_7;
input 	cfg_twr_wire_0;
input 	cfg_twr_wire_1;
input 	cfg_twr_wire_2;
input 	cfg_twr_wire_3;
input 	afi_mem_clk_disable_0;
input 	cfg_dramconfig_wire_0;
input 	cfg_dramconfig_wire_1;
input 	cfg_dramconfig_wire_2;
input 	cfg_dramconfig_wire_3;
input 	cfg_dramconfig_wire_4;
input 	cfg_dramconfig_wire_5;
input 	cfg_dramconfig_wire_6;
input 	cfg_dramconfig_wire_7;
input 	cfg_dramconfig_wire_8;
input 	cfg_dramconfig_wire_9;
input 	cfg_dramconfig_wire_10;
input 	cfg_dramconfig_wire_11;
input 	cfg_dramconfig_wire_12;
input 	cfg_dramconfig_wire_13;
input 	cfg_dramconfig_wire_14;
input 	cfg_dramconfig_wire_15;
input 	cfg_dramconfig_wire_16;
input 	cfg_dramconfig_wire_17;
input 	cfg_dramconfig_wire_18;
input 	cfg_dramconfig_wire_19;
input 	cfg_dramconfig_wire_20;
output 	ctl_clk;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_hps_sdram_p0_acv_hard_memphy umemphy(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.afi_cal_fail(afi_cal_fail),
	.afi_cal_success(afi_cal_success),
	.afi_rdata_valid({afi_rdata_valid_0}),
	.ctl_reset_n(ctl_reset_n),
	.afi_rdata({afi_rdata_79,afi_rdata_78,afi_rdata_77,afi_rdata_76,afi_rdata_75,afi_rdata_74,afi_rdata_73,afi_rdata_72,afi_rdata_71,afi_rdata_70,afi_rdata_69,afi_rdata_68,afi_rdata_67,afi_rdata_66,afi_rdata_65,afi_rdata_64,afi_rdata_63,afi_rdata_62,afi_rdata_61,afi_rdata_60,afi_rdata_59,
afi_rdata_58,afi_rdata_57,afi_rdata_56,afi_rdata_55,afi_rdata_54,afi_rdata_53,afi_rdata_52,afi_rdata_51,afi_rdata_50,afi_rdata_49,afi_rdata_48,afi_rdata_47,afi_rdata_46,afi_rdata_45,afi_rdata_44,afi_rdata_43,afi_rdata_42,afi_rdata_41,afi_rdata_40,afi_rdata_39,afi_rdata_38,
afi_rdata_37,afi_rdata_36,afi_rdata_35,afi_rdata_34,afi_rdata_33,afi_rdata_32,afi_rdata_31,afi_rdata_30,afi_rdata_29,afi_rdata_28,afi_rdata_27,afi_rdata_26,afi_rdata_25,afi_rdata_24,afi_rdata_23,afi_rdata_22,afi_rdata_21,afi_rdata_20,afi_rdata_19,afi_rdata_18,afi_rdata_17,
afi_rdata_16,afi_rdata_15,afi_rdata_14,afi_rdata_13,afi_rdata_12,afi_rdata_11,afi_rdata_10,afi_rdata_9,afi_rdata_8,afi_rdata_7,afi_rdata_6,afi_rdata_5,afi_rdata_4,afi_rdata_3,afi_rdata_2,afi_rdata_1,afi_rdata_0}),
	.afi_wlat({afi_wlat_3,afi_wlat_2,afi_wlat_1,afi_wlat_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.afi_cas_n({afi_cas_n_0}),
	.afi_ras_n({afi_ras_n_0}),
	.afi_rst_n({afi_rst_n_0}),
	.afi_we_n({afi_we_n_0}),
	.afi_addr({afi_addr_19,afi_addr_18,afi_addr_17,afi_addr_16,afi_addr_15,afi_addr_14,afi_addr_13,afi_addr_12,afi_addr_11,afi_addr_10,afi_addr_9,afi_addr_8,afi_addr_7,afi_addr_6,afi_addr_5,afi_addr_4,afi_addr_3,afi_addr_2,afi_addr_1,afi_addr_0}),
	.afi_ba({afi_ba_2,afi_ba_1,afi_ba_0}),
	.afi_cke({afi_cke_1,afi_cke_0}),
	.afi_cs_n({afi_cs_n_1,afi_cs_n_0}),
	.afi_dm({afi_dm_int_9,afi_dm_int_8,afi_dm_int_7,afi_dm_int_6,afi_dm_int_5,afi_dm_int_4,afi_dm_int_3,afi_dm_int_2,afi_dm_int_1,afi_dm_int_0}),
	.afi_dqs_burst({afi_dqs_burst_4,afi_dqs_burst_3,afi_dqs_burst_2,afi_dqs_burst_1,afi_dqs_burst_0}),
	.afi_odt({afi_odt_1,afi_odt_0}),
	.afi_rdata_en({afi_rdata_en_4,afi_rdata_en_3,afi_rdata_en_2,afi_rdata_en_1,afi_rdata_en_0}),
	.afi_rdata_en_full({afi_rdata_en_full_4,afi_rdata_en_full_3,afi_rdata_en_full_2,afi_rdata_en_full_1,afi_rdata_en_full_0}),
	.afi_wdata({afi_wdata_int_79,afi_wdata_int_78,afi_wdata_int_77,afi_wdata_int_76,afi_wdata_int_75,afi_wdata_int_74,afi_wdata_int_73,afi_wdata_int_72,afi_wdata_int_71,afi_wdata_int_70,afi_wdata_int_69,afi_wdata_int_68,afi_wdata_int_67,afi_wdata_int_66,afi_wdata_int_65,afi_wdata_int_64,
afi_wdata_int_63,afi_wdata_int_62,afi_wdata_int_61,afi_wdata_int_60,afi_wdata_int_59,afi_wdata_int_58,afi_wdata_int_57,afi_wdata_int_56,afi_wdata_int_55,afi_wdata_int_54,afi_wdata_int_53,afi_wdata_int_52,afi_wdata_int_51,afi_wdata_int_50,afi_wdata_int_49,afi_wdata_int_48,
afi_wdata_int_47,afi_wdata_int_46,afi_wdata_int_45,afi_wdata_int_44,afi_wdata_int_43,afi_wdata_int_42,afi_wdata_int_41,afi_wdata_int_40,afi_wdata_int_39,afi_wdata_int_38,afi_wdata_int_37,afi_wdata_int_36,afi_wdata_int_35,afi_wdata_int_34,afi_wdata_int_33,afi_wdata_int_32,
afi_wdata_int_31,afi_wdata_int_30,afi_wdata_int_29,afi_wdata_int_28,afi_wdata_int_27,afi_wdata_int_26,afi_wdata_int_25,afi_wdata_int_24,afi_wdata_int_23,afi_wdata_int_22,afi_wdata_int_21,afi_wdata_int_20,afi_wdata_int_19,afi_wdata_int_18,afi_wdata_int_17,afi_wdata_int_16,
afi_wdata_int_15,afi_wdata_int_14,afi_wdata_int_13,afi_wdata_int_12,afi_wdata_int_11,afi_wdata_int_10,afi_wdata_int_9,afi_wdata_int_8,afi_wdata_int_7,afi_wdata_int_6,afi_wdata_int_5,afi_wdata_int_4,afi_wdata_int_3,afi_wdata_int_2,afi_wdata_int_1,afi_wdata_int_0}),
	.afi_wdata_valid({afi_wdata_valid_4,afi_wdata_valid_3,afi_wdata_valid_2,afi_wdata_valid_1,afi_wdata_valid_0}),
	.cfg_addlat({gnd,gnd,gnd,cfg_addlat_wire_4,cfg_addlat_wire_3,cfg_addlat_wire_2,cfg_addlat_wire_1,cfg_addlat_wire_0}),
	.cfg_bankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth_wire_2,cfg_bankaddrwidth_wire_1,cfg_bankaddrwidth_wire_0}),
	.cfg_caswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat_wire_3,cfg_caswrlat_wire_2,cfg_caswrlat_wire_1,cfg_caswrlat_wire_0}),
	.cfg_coladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth_wire_4,cfg_coladdrwidth_wire_3,cfg_coladdrwidth_wire_2,cfg_coladdrwidth_wire_1,cfg_coladdrwidth_wire_0}),
	.cfg_csaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth_wire_2,cfg_csaddrwidth_wire_1,cfg_csaddrwidth_wire_0}),
	.cfg_devicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth_wire_3,cfg_devicewidth_wire_2,cfg_devicewidth_wire_1,cfg_devicewidth_wire_0}),
	.cfg_interfacewidth({cfg_interfacewidth_wire_7,cfg_interfacewidth_wire_6,cfg_interfacewidth_wire_5,cfg_interfacewidth_wire_4,cfg_interfacewidth_wire_3,cfg_interfacewidth_wire_2,cfg_interfacewidth_wire_1,cfg_interfacewidth_wire_0}),
	.cfg_rowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth_wire_4,cfg_rowaddrwidth_wire_3,cfg_rowaddrwidth_wire_2,cfg_rowaddrwidth_wire_1,cfg_rowaddrwidth_wire_0}),
	.cfg_tcl({gnd,gnd,gnd,cfg_tcl_wire_4,cfg_tcl_wire_3,cfg_tcl_wire_2,cfg_tcl_wire_1,cfg_tcl_wire_0}),
	.cfg_tmrd({gnd,gnd,gnd,gnd,cfg_tmrd_wire_3,cfg_tmrd_wire_2,cfg_tmrd_wire_1,cfg_tmrd_wire_0}),
	.cfg_trefi({gnd,gnd,gnd,cfg_trefi_wire_12,cfg_trefi_wire_11,cfg_trefi_wire_10,cfg_trefi_wire_9,cfg_trefi_wire_8,cfg_trefi_wire_7,cfg_trefi_wire_6,cfg_trefi_wire_5,cfg_trefi_wire_4,cfg_trefi_wire_3,cfg_trefi_wire_2,cfg_trefi_wire_1,cfg_trefi_wire_0}),
	.cfg_trfc({cfg_trfc_wire_7,cfg_trfc_wire_6,cfg_trfc_wire_5,cfg_trfc_wire_4,cfg_trfc_wire_3,cfg_trfc_wire_2,cfg_trfc_wire_1,cfg_trfc_wire_0}),
	.cfg_twr({gnd,gnd,gnd,gnd,cfg_twr_wire_3,cfg_twr_wire_2,cfg_twr_wire_1,cfg_twr_wire_0}),
	.afi_mem_clk_disable({afi_mem_clk_disable_0}),
	.cfg_dramconfig({gnd,gnd,gnd,cfg_dramconfig_wire_20,cfg_dramconfig_wire_19,cfg_dramconfig_wire_18,cfg_dramconfig_wire_17,cfg_dramconfig_wire_16,cfg_dramconfig_wire_15,cfg_dramconfig_wire_14,cfg_dramconfig_wire_13,cfg_dramconfig_wire_12,cfg_dramconfig_wire_11,cfg_dramconfig_wire_10,
cfg_dramconfig_wire_9,cfg_dramconfig_wire_8,cfg_dramconfig_wire_7,cfg_dramconfig_wire_6,cfg_dramconfig_wire_5,cfg_dramconfig_wire_4,cfg_dramconfig_wire_3,cfg_dramconfig_wire_2,cfg_dramconfig_wire_1,cfg_dramconfig_wire_0}),
	.ctl_clk(ctl_clk),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module terminal_qsys_hps_sdram_p0_acv_hard_memphy (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	afi_cal_fail,
	afi_cal_success,
	afi_rdata_valid,
	ctl_reset_n,
	afi_rdata,
	afi_wlat,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	afi_cas_n,
	afi_ras_n,
	afi_rst_n,
	afi_we_n,
	afi_addr,
	afi_ba,
	afi_cke,
	afi_cs_n,
	afi_dm,
	afi_dqs_burst,
	afi_odt,
	afi_rdata_en,
	afi_rdata_en_full,
	afi_wdata,
	afi_wdata_valid,
	cfg_addlat,
	cfg_bankaddrwidth,
	cfg_caswrlat,
	cfg_coladdrwidth,
	cfg_csaddrwidth,
	cfg_devicewidth,
	cfg_interfacewidth,
	cfg_rowaddrwidth,
	cfg_tcl,
	cfg_tmrd,
	cfg_trefi,
	cfg_trfc,
	cfg_twr,
	afi_mem_clk_disable,
	cfg_dramconfig,
	ctl_clk,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
output 	afi_cal_fail;
output 	afi_cal_success;
output 	[0:0] afi_rdata_valid;
output 	ctl_reset_n;
output 	[79:0] afi_rdata;
output 	[3:0] afi_wlat;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
input 	[0:0] afi_cas_n;
input 	[0:0] afi_ras_n;
input 	[0:0] afi_rst_n;
input 	[0:0] afi_we_n;
input 	[19:0] afi_addr;
input 	[2:0] afi_ba;
input 	[1:0] afi_cke;
input 	[1:0] afi_cs_n;
input 	[9:0] afi_dm;
input 	[4:0] afi_dqs_burst;
input 	[1:0] afi_odt;
input 	[4:0] afi_rdata_en;
input 	[4:0] afi_rdata_en_full;
input 	[79:0] afi_wdata;
input 	[4:0] afi_wdata_valid;
input 	[7:0] cfg_addlat;
input 	[7:0] cfg_bankaddrwidth;
input 	[7:0] cfg_caswrlat;
input 	[7:0] cfg_coladdrwidth;
input 	[7:0] cfg_csaddrwidth;
input 	[7:0] cfg_devicewidth;
input 	[7:0] cfg_interfacewidth;
input 	[7:0] cfg_rowaddrwidth;
input 	[7:0] cfg_tcl;
input 	[7:0] cfg_tmrd;
input 	[15:0] cfg_trefi;
input 	[7:0] cfg_trfc;
input 	[7:0] cfg_twr;
input 	[0:0] afi_mem_clk_disable;
input 	[23:0] cfg_dramconfig;
output 	ctl_clk;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \memphy_ldc|leveled_hr_clocks[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ;
wire \uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ;
wire \phy_ddio_address[0] ;
wire \phy_ddio_address[1] ;
wire \phy_ddio_address[2] ;
wire \phy_ddio_address[3] ;
wire \phy_ddio_address[4] ;
wire \phy_ddio_address[5] ;
wire \phy_ddio_address[6] ;
wire \phy_ddio_address[7] ;
wire \phy_ddio_address[8] ;
wire \phy_ddio_address[9] ;
wire \phy_ddio_address[10] ;
wire \phy_ddio_address[11] ;
wire \phy_ddio_address[12] ;
wire \phy_ddio_address[13] ;
wire \phy_ddio_address[14] ;
wire \phy_ddio_address[15] ;
wire \phy_ddio_address[16] ;
wire \phy_ddio_address[17] ;
wire \phy_ddio_address[18] ;
wire \phy_ddio_address[19] ;
wire \phy_ddio_address[20] ;
wire \phy_ddio_address[21] ;
wire \phy_ddio_address[22] ;
wire \phy_ddio_address[23] ;
wire \phy_ddio_address[24] ;
wire \phy_ddio_address[25] ;
wire \phy_ddio_address[26] ;
wire \phy_ddio_address[27] ;
wire \phy_ddio_address[28] ;
wire \phy_ddio_address[29] ;
wire \phy_ddio_address[30] ;
wire \phy_ddio_address[31] ;
wire \phy_ddio_address[32] ;
wire \phy_ddio_address[33] ;
wire \phy_ddio_address[34] ;
wire \phy_ddio_address[35] ;
wire \phy_ddio_address[36] ;
wire \phy_ddio_address[37] ;
wire \phy_ddio_address[38] ;
wire \phy_ddio_address[39] ;
wire \phy_ddio_address[40] ;
wire \phy_ddio_address[41] ;
wire \phy_ddio_address[42] ;
wire \phy_ddio_address[43] ;
wire \phy_ddio_address[44] ;
wire \phy_ddio_address[45] ;
wire \phy_ddio_address[46] ;
wire \phy_ddio_address[47] ;
wire \phy_ddio_address[48] ;
wire \phy_ddio_address[49] ;
wire \phy_ddio_address[50] ;
wire \phy_ddio_address[51] ;
wire \phy_ddio_address[52] ;
wire \phy_ddio_address[53] ;
wire \phy_ddio_address[54] ;
wire \phy_ddio_address[55] ;
wire \phy_ddio_address[56] ;
wire \phy_ddio_address[57] ;
wire \phy_ddio_address[58] ;
wire \phy_ddio_address[59] ;
wire \phy_ddio_bank[0] ;
wire \phy_ddio_bank[1] ;
wire \phy_ddio_bank[2] ;
wire \phy_ddio_bank[3] ;
wire \phy_ddio_bank[4] ;
wire \phy_ddio_bank[5] ;
wire \phy_ddio_bank[6] ;
wire \phy_ddio_bank[7] ;
wire \phy_ddio_bank[8] ;
wire \phy_ddio_bank[9] ;
wire \phy_ddio_bank[10] ;
wire \phy_ddio_bank[11] ;
wire \phy_ddio_cas_n[0] ;
wire \phy_ddio_cas_n[1] ;
wire \phy_ddio_cas_n[2] ;
wire \phy_ddio_cas_n[3] ;
wire \phy_ddio_ck[0] ;
wire \phy_ddio_ck[1] ;
wire \phy_ddio_cke[0] ;
wire \phy_ddio_cke[1] ;
wire \phy_ddio_cke[2] ;
wire \phy_ddio_cke[3] ;
wire \phy_ddio_cs_n[0] ;
wire \phy_ddio_cs_n[1] ;
wire \phy_ddio_cs_n[2] ;
wire \phy_ddio_cs_n[3] ;
wire \phy_ddio_dmdout[0] ;
wire \phy_ddio_dmdout[1] ;
wire \phy_ddio_dmdout[2] ;
wire \phy_ddio_dmdout[3] ;
wire \phy_ddio_dmdout[4] ;
wire \phy_ddio_dmdout[5] ;
wire \phy_ddio_dmdout[6] ;
wire \phy_ddio_dmdout[7] ;
wire \phy_ddio_dmdout[8] ;
wire \phy_ddio_dmdout[9] ;
wire \phy_ddio_dmdout[10] ;
wire \phy_ddio_dmdout[11] ;
wire \phy_ddio_dmdout[12] ;
wire \phy_ddio_dmdout[13] ;
wire \phy_ddio_dmdout[14] ;
wire \phy_ddio_dmdout[15] ;
wire \phy_ddio_dqdout[0] ;
wire \phy_ddio_dqdout[1] ;
wire \phy_ddio_dqdout[2] ;
wire \phy_ddio_dqdout[3] ;
wire \phy_ddio_dqdout[4] ;
wire \phy_ddio_dqdout[5] ;
wire \phy_ddio_dqdout[6] ;
wire \phy_ddio_dqdout[7] ;
wire \phy_ddio_dqdout[8] ;
wire \phy_ddio_dqdout[9] ;
wire \phy_ddio_dqdout[10] ;
wire \phy_ddio_dqdout[11] ;
wire \phy_ddio_dqdout[12] ;
wire \phy_ddio_dqdout[13] ;
wire \phy_ddio_dqdout[14] ;
wire \phy_ddio_dqdout[15] ;
wire \phy_ddio_dqdout[16] ;
wire \phy_ddio_dqdout[17] ;
wire \phy_ddio_dqdout[18] ;
wire \phy_ddio_dqdout[19] ;
wire \phy_ddio_dqdout[20] ;
wire \phy_ddio_dqdout[21] ;
wire \phy_ddio_dqdout[22] ;
wire \phy_ddio_dqdout[23] ;
wire \phy_ddio_dqdout[24] ;
wire \phy_ddio_dqdout[25] ;
wire \phy_ddio_dqdout[26] ;
wire \phy_ddio_dqdout[27] ;
wire \phy_ddio_dqdout[28] ;
wire \phy_ddio_dqdout[29] ;
wire \phy_ddio_dqdout[30] ;
wire \phy_ddio_dqdout[31] ;
wire \phy_ddio_dqdout[36] ;
wire \phy_ddio_dqdout[37] ;
wire \phy_ddio_dqdout[38] ;
wire \phy_ddio_dqdout[39] ;
wire \phy_ddio_dqdout[40] ;
wire \phy_ddio_dqdout[41] ;
wire \phy_ddio_dqdout[42] ;
wire \phy_ddio_dqdout[43] ;
wire \phy_ddio_dqdout[44] ;
wire \phy_ddio_dqdout[45] ;
wire \phy_ddio_dqdout[46] ;
wire \phy_ddio_dqdout[47] ;
wire \phy_ddio_dqdout[48] ;
wire \phy_ddio_dqdout[49] ;
wire \phy_ddio_dqdout[50] ;
wire \phy_ddio_dqdout[51] ;
wire \phy_ddio_dqdout[52] ;
wire \phy_ddio_dqdout[53] ;
wire \phy_ddio_dqdout[54] ;
wire \phy_ddio_dqdout[55] ;
wire \phy_ddio_dqdout[56] ;
wire \phy_ddio_dqdout[57] ;
wire \phy_ddio_dqdout[58] ;
wire \phy_ddio_dqdout[59] ;
wire \phy_ddio_dqdout[60] ;
wire \phy_ddio_dqdout[61] ;
wire \phy_ddio_dqdout[62] ;
wire \phy_ddio_dqdout[63] ;
wire \phy_ddio_dqdout[64] ;
wire \phy_ddio_dqdout[65] ;
wire \phy_ddio_dqdout[66] ;
wire \phy_ddio_dqdout[67] ;
wire \phy_ddio_dqdout[72] ;
wire \phy_ddio_dqdout[73] ;
wire \phy_ddio_dqdout[74] ;
wire \phy_ddio_dqdout[75] ;
wire \phy_ddio_dqdout[76] ;
wire \phy_ddio_dqdout[77] ;
wire \phy_ddio_dqdout[78] ;
wire \phy_ddio_dqdout[79] ;
wire \phy_ddio_dqdout[80] ;
wire \phy_ddio_dqdout[81] ;
wire \phy_ddio_dqdout[82] ;
wire \phy_ddio_dqdout[83] ;
wire \phy_ddio_dqdout[84] ;
wire \phy_ddio_dqdout[85] ;
wire \phy_ddio_dqdout[86] ;
wire \phy_ddio_dqdout[87] ;
wire \phy_ddio_dqdout[88] ;
wire \phy_ddio_dqdout[89] ;
wire \phy_ddio_dqdout[90] ;
wire \phy_ddio_dqdout[91] ;
wire \phy_ddio_dqdout[92] ;
wire \phy_ddio_dqdout[93] ;
wire \phy_ddio_dqdout[94] ;
wire \phy_ddio_dqdout[95] ;
wire \phy_ddio_dqdout[96] ;
wire \phy_ddio_dqdout[97] ;
wire \phy_ddio_dqdout[98] ;
wire \phy_ddio_dqdout[99] ;
wire \phy_ddio_dqdout[100] ;
wire \phy_ddio_dqdout[101] ;
wire \phy_ddio_dqdout[102] ;
wire \phy_ddio_dqdout[103] ;
wire \phy_ddio_dqdout[108] ;
wire \phy_ddio_dqdout[109] ;
wire \phy_ddio_dqdout[110] ;
wire \phy_ddio_dqdout[111] ;
wire \phy_ddio_dqdout[112] ;
wire \phy_ddio_dqdout[113] ;
wire \phy_ddio_dqdout[114] ;
wire \phy_ddio_dqdout[115] ;
wire \phy_ddio_dqdout[116] ;
wire \phy_ddio_dqdout[117] ;
wire \phy_ddio_dqdout[118] ;
wire \phy_ddio_dqdout[119] ;
wire \phy_ddio_dqdout[120] ;
wire \phy_ddio_dqdout[121] ;
wire \phy_ddio_dqdout[122] ;
wire \phy_ddio_dqdout[123] ;
wire \phy_ddio_dqdout[124] ;
wire \phy_ddio_dqdout[125] ;
wire \phy_ddio_dqdout[126] ;
wire \phy_ddio_dqdout[127] ;
wire \phy_ddio_dqdout[128] ;
wire \phy_ddio_dqdout[129] ;
wire \phy_ddio_dqdout[130] ;
wire \phy_ddio_dqdout[131] ;
wire \phy_ddio_dqdout[132] ;
wire \phy_ddio_dqdout[133] ;
wire \phy_ddio_dqdout[134] ;
wire \phy_ddio_dqdout[135] ;
wire \phy_ddio_dqdout[136] ;
wire \phy_ddio_dqdout[137] ;
wire \phy_ddio_dqdout[138] ;
wire \phy_ddio_dqdout[139] ;
wire \phy_ddio_dqoe[0] ;
wire \phy_ddio_dqoe[1] ;
wire \phy_ddio_dqoe[2] ;
wire \phy_ddio_dqoe[3] ;
wire \phy_ddio_dqoe[4] ;
wire \phy_ddio_dqoe[5] ;
wire \phy_ddio_dqoe[6] ;
wire \phy_ddio_dqoe[7] ;
wire \phy_ddio_dqoe[8] ;
wire \phy_ddio_dqoe[9] ;
wire \phy_ddio_dqoe[10] ;
wire \phy_ddio_dqoe[11] ;
wire \phy_ddio_dqoe[12] ;
wire \phy_ddio_dqoe[13] ;
wire \phy_ddio_dqoe[14] ;
wire \phy_ddio_dqoe[15] ;
wire \phy_ddio_dqoe[18] ;
wire \phy_ddio_dqoe[19] ;
wire \phy_ddio_dqoe[20] ;
wire \phy_ddio_dqoe[21] ;
wire \phy_ddio_dqoe[22] ;
wire \phy_ddio_dqoe[23] ;
wire \phy_ddio_dqoe[24] ;
wire \phy_ddio_dqoe[25] ;
wire \phy_ddio_dqoe[26] ;
wire \phy_ddio_dqoe[27] ;
wire \phy_ddio_dqoe[28] ;
wire \phy_ddio_dqoe[29] ;
wire \phy_ddio_dqoe[30] ;
wire \phy_ddio_dqoe[31] ;
wire \phy_ddio_dqoe[32] ;
wire \phy_ddio_dqoe[33] ;
wire \phy_ddio_dqoe[36] ;
wire \phy_ddio_dqoe[37] ;
wire \phy_ddio_dqoe[38] ;
wire \phy_ddio_dqoe[39] ;
wire \phy_ddio_dqoe[40] ;
wire \phy_ddio_dqoe[41] ;
wire \phy_ddio_dqoe[42] ;
wire \phy_ddio_dqoe[43] ;
wire \phy_ddio_dqoe[44] ;
wire \phy_ddio_dqoe[45] ;
wire \phy_ddio_dqoe[46] ;
wire \phy_ddio_dqoe[47] ;
wire \phy_ddio_dqoe[48] ;
wire \phy_ddio_dqoe[49] ;
wire \phy_ddio_dqoe[50] ;
wire \phy_ddio_dqoe[51] ;
wire \phy_ddio_dqoe[54] ;
wire \phy_ddio_dqoe[55] ;
wire \phy_ddio_dqoe[56] ;
wire \phy_ddio_dqoe[57] ;
wire \phy_ddio_dqoe[58] ;
wire \phy_ddio_dqoe[59] ;
wire \phy_ddio_dqoe[60] ;
wire \phy_ddio_dqoe[61] ;
wire \phy_ddio_dqoe[62] ;
wire \phy_ddio_dqoe[63] ;
wire \phy_ddio_dqoe[64] ;
wire \phy_ddio_dqoe[65] ;
wire \phy_ddio_dqoe[66] ;
wire \phy_ddio_dqoe[67] ;
wire \phy_ddio_dqoe[68] ;
wire \phy_ddio_dqoe[69] ;
wire \phy_ddio_dqs_dout[0] ;
wire \phy_ddio_dqs_dout[1] ;
wire \phy_ddio_dqs_dout[2] ;
wire \phy_ddio_dqs_dout[3] ;
wire \phy_ddio_dqs_dout[4] ;
wire \phy_ddio_dqs_dout[5] ;
wire \phy_ddio_dqs_dout[6] ;
wire \phy_ddio_dqs_dout[7] ;
wire \phy_ddio_dqs_dout[8] ;
wire \phy_ddio_dqs_dout[9] ;
wire \phy_ddio_dqs_dout[10] ;
wire \phy_ddio_dqs_dout[11] ;
wire \phy_ddio_dqs_dout[12] ;
wire \phy_ddio_dqs_dout[13] ;
wire \phy_ddio_dqs_dout[14] ;
wire \phy_ddio_dqs_dout[15] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[0] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[1] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[2] ;
wire \phy_ddio_dqslogic_aclr_fifoctrl[3] ;
wire \phy_ddio_dqslogic_aclr_pstamble[0] ;
wire \phy_ddio_dqslogic_aclr_pstamble[1] ;
wire \phy_ddio_dqslogic_aclr_pstamble[2] ;
wire \phy_ddio_dqslogic_aclr_pstamble[3] ;
wire \phy_ddio_dqslogic_dqsena[0] ;
wire \phy_ddio_dqslogic_dqsena[1] ;
wire \phy_ddio_dqslogic_dqsena[2] ;
wire \phy_ddio_dqslogic_dqsena[3] ;
wire \phy_ddio_dqslogic_dqsena[4] ;
wire \phy_ddio_dqslogic_dqsena[5] ;
wire \phy_ddio_dqslogic_dqsena[6] ;
wire \phy_ddio_dqslogic_dqsena[7] ;
wire \phy_ddio_dqslogic_fiforeset[0] ;
wire \phy_ddio_dqslogic_fiforeset[1] ;
wire \phy_ddio_dqslogic_fiforeset[2] ;
wire \phy_ddio_dqslogic_fiforeset[3] ;
wire \phy_ddio_dqslogic_incrdataen[0] ;
wire \phy_ddio_dqslogic_incrdataen[1] ;
wire \phy_ddio_dqslogic_incrdataen[2] ;
wire \phy_ddio_dqslogic_incrdataen[3] ;
wire \phy_ddio_dqslogic_incrdataen[4] ;
wire \phy_ddio_dqslogic_incrdataen[5] ;
wire \phy_ddio_dqslogic_incrdataen[6] ;
wire \phy_ddio_dqslogic_incrdataen[7] ;
wire \phy_ddio_dqslogic_incwrptr[0] ;
wire \phy_ddio_dqslogic_incwrptr[1] ;
wire \phy_ddio_dqslogic_incwrptr[2] ;
wire \phy_ddio_dqslogic_incwrptr[3] ;
wire \phy_ddio_dqslogic_incwrptr[4] ;
wire \phy_ddio_dqslogic_incwrptr[5] ;
wire \phy_ddio_dqslogic_incwrptr[6] ;
wire \phy_ddio_dqslogic_incwrptr[7] ;
wire \phy_ddio_dqslogic_oct[0] ;
wire \phy_ddio_dqslogic_oct[1] ;
wire \phy_ddio_dqslogic_oct[2] ;
wire \phy_ddio_dqslogic_oct[3] ;
wire \phy_ddio_dqslogic_oct[4] ;
wire \phy_ddio_dqslogic_oct[5] ;
wire \phy_ddio_dqslogic_oct[6] ;
wire \phy_ddio_dqslogic_oct[7] ;
wire \phy_ddio_dqslogic_readlatency[0] ;
wire \phy_ddio_dqslogic_readlatency[1] ;
wire \phy_ddio_dqslogic_readlatency[2] ;
wire \phy_ddio_dqslogic_readlatency[3] ;
wire \phy_ddio_dqslogic_readlatency[4] ;
wire \phy_ddio_dqslogic_readlatency[5] ;
wire \phy_ddio_dqslogic_readlatency[6] ;
wire \phy_ddio_dqslogic_readlatency[7] ;
wire \phy_ddio_dqslogic_readlatency[8] ;
wire \phy_ddio_dqslogic_readlatency[9] ;
wire \phy_ddio_dqslogic_readlatency[10] ;
wire \phy_ddio_dqslogic_readlatency[11] ;
wire \phy_ddio_dqslogic_readlatency[12] ;
wire \phy_ddio_dqslogic_readlatency[13] ;
wire \phy_ddio_dqslogic_readlatency[14] ;
wire \phy_ddio_dqslogic_readlatency[15] ;
wire \phy_ddio_dqslogic_readlatency[16] ;
wire \phy_ddio_dqslogic_readlatency[17] ;
wire \phy_ddio_dqslogic_readlatency[18] ;
wire \phy_ddio_dqslogic_readlatency[19] ;
wire \phy_ddio_dqs_oe[0] ;
wire \phy_ddio_dqs_oe[1] ;
wire \phy_ddio_dqs_oe[2] ;
wire \phy_ddio_dqs_oe[3] ;
wire \phy_ddio_dqs_oe[4] ;
wire \phy_ddio_dqs_oe[5] ;
wire \phy_ddio_dqs_oe[6] ;
wire \phy_ddio_dqs_oe[7] ;
wire \phy_ddio_odt[0] ;
wire \phy_ddio_odt[1] ;
wire \phy_ddio_odt[2] ;
wire \phy_ddio_odt[3] ;
wire \phy_ddio_ras_n[0] ;
wire \phy_ddio_ras_n[1] ;
wire \phy_ddio_ras_n[2] ;
wire \phy_ddio_ras_n[3] ;
wire \phy_ddio_reset_n[0] ;
wire \phy_ddio_reset_n[1] ;
wire \phy_ddio_reset_n[2] ;
wire \phy_ddio_reset_n[3] ;
wire \phy_ddio_we_n[0] ;
wire \phy_ddio_we_n[1] ;
wire \phy_ddio_we_n[2] ;
wire \phy_ddio_we_n[3] ;

wire [79:0] hphy_inst_AFIRDATA_bus;
wire [3:0] hphy_inst_AFIWLAT_bus;
wire [63:0] hphy_inst_PHYDDIOADDRDOUT_bus;
wire [11:0] hphy_inst_PHYDDIOBADOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOCKDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCKEDOUT_bus;
wire [7:0] hphy_inst_PHYDDIOCSNDOUT_bus;
wire [19:0] hphy_inst_PHYDDIODMDOUT_bus;
wire [179:0] hphy_inst_PHYDDIODQDOUT_bus;
wire [89:0] hphy_inst_PHYDDIODQOE_bus;
wire [19:0] hphy_inst_PHYDDIODQSDOUT_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICDQSENA_bus;
wire [4:0] hphy_inst_PHYDDIODQSLOGICFIFORESET_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus;
wire [9:0] hphy_inst_PHYDDIODQSLOGICOCT_bus;
wire [24:0] hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus;
wire [9:0] hphy_inst_PHYDDIODQSOE_bus;
wire [7:0] hphy_inst_PHYDDIOODTDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORASNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIORESETNDOUT_bus;
wire [3:0] hphy_inst_PHYDDIOWENDOUT_bus;

assign afi_rdata[0] = hphy_inst_AFIRDATA_bus[0];
assign afi_rdata[1] = hphy_inst_AFIRDATA_bus[1];
assign afi_rdata[2] = hphy_inst_AFIRDATA_bus[2];
assign afi_rdata[3] = hphy_inst_AFIRDATA_bus[3];
assign afi_rdata[4] = hphy_inst_AFIRDATA_bus[4];
assign afi_rdata[5] = hphy_inst_AFIRDATA_bus[5];
assign afi_rdata[6] = hphy_inst_AFIRDATA_bus[6];
assign afi_rdata[7] = hphy_inst_AFIRDATA_bus[7];
assign afi_rdata[8] = hphy_inst_AFIRDATA_bus[8];
assign afi_rdata[9] = hphy_inst_AFIRDATA_bus[9];
assign afi_rdata[10] = hphy_inst_AFIRDATA_bus[10];
assign afi_rdata[11] = hphy_inst_AFIRDATA_bus[11];
assign afi_rdata[12] = hphy_inst_AFIRDATA_bus[12];
assign afi_rdata[13] = hphy_inst_AFIRDATA_bus[13];
assign afi_rdata[14] = hphy_inst_AFIRDATA_bus[14];
assign afi_rdata[15] = hphy_inst_AFIRDATA_bus[15];
assign afi_rdata[16] = hphy_inst_AFIRDATA_bus[16];
assign afi_rdata[17] = hphy_inst_AFIRDATA_bus[17];
assign afi_rdata[18] = hphy_inst_AFIRDATA_bus[18];
assign afi_rdata[19] = hphy_inst_AFIRDATA_bus[19];
assign afi_rdata[20] = hphy_inst_AFIRDATA_bus[20];
assign afi_rdata[21] = hphy_inst_AFIRDATA_bus[21];
assign afi_rdata[22] = hphy_inst_AFIRDATA_bus[22];
assign afi_rdata[23] = hphy_inst_AFIRDATA_bus[23];
assign afi_rdata[24] = hphy_inst_AFIRDATA_bus[24];
assign afi_rdata[25] = hphy_inst_AFIRDATA_bus[25];
assign afi_rdata[26] = hphy_inst_AFIRDATA_bus[26];
assign afi_rdata[27] = hphy_inst_AFIRDATA_bus[27];
assign afi_rdata[28] = hphy_inst_AFIRDATA_bus[28];
assign afi_rdata[29] = hphy_inst_AFIRDATA_bus[29];
assign afi_rdata[30] = hphy_inst_AFIRDATA_bus[30];
assign afi_rdata[31] = hphy_inst_AFIRDATA_bus[31];
assign afi_rdata[32] = hphy_inst_AFIRDATA_bus[32];
assign afi_rdata[33] = hphy_inst_AFIRDATA_bus[33];
assign afi_rdata[34] = hphy_inst_AFIRDATA_bus[34];
assign afi_rdata[35] = hphy_inst_AFIRDATA_bus[35];
assign afi_rdata[36] = hphy_inst_AFIRDATA_bus[36];
assign afi_rdata[37] = hphy_inst_AFIRDATA_bus[37];
assign afi_rdata[38] = hphy_inst_AFIRDATA_bus[38];
assign afi_rdata[39] = hphy_inst_AFIRDATA_bus[39];
assign afi_rdata[40] = hphy_inst_AFIRDATA_bus[40];
assign afi_rdata[41] = hphy_inst_AFIRDATA_bus[41];
assign afi_rdata[42] = hphy_inst_AFIRDATA_bus[42];
assign afi_rdata[43] = hphy_inst_AFIRDATA_bus[43];
assign afi_rdata[44] = hphy_inst_AFIRDATA_bus[44];
assign afi_rdata[45] = hphy_inst_AFIRDATA_bus[45];
assign afi_rdata[46] = hphy_inst_AFIRDATA_bus[46];
assign afi_rdata[47] = hphy_inst_AFIRDATA_bus[47];
assign afi_rdata[48] = hphy_inst_AFIRDATA_bus[48];
assign afi_rdata[49] = hphy_inst_AFIRDATA_bus[49];
assign afi_rdata[50] = hphy_inst_AFIRDATA_bus[50];
assign afi_rdata[51] = hphy_inst_AFIRDATA_bus[51];
assign afi_rdata[52] = hphy_inst_AFIRDATA_bus[52];
assign afi_rdata[53] = hphy_inst_AFIRDATA_bus[53];
assign afi_rdata[54] = hphy_inst_AFIRDATA_bus[54];
assign afi_rdata[55] = hphy_inst_AFIRDATA_bus[55];
assign afi_rdata[56] = hphy_inst_AFIRDATA_bus[56];
assign afi_rdata[57] = hphy_inst_AFIRDATA_bus[57];
assign afi_rdata[58] = hphy_inst_AFIRDATA_bus[58];
assign afi_rdata[59] = hphy_inst_AFIRDATA_bus[59];
assign afi_rdata[60] = hphy_inst_AFIRDATA_bus[60];
assign afi_rdata[61] = hphy_inst_AFIRDATA_bus[61];
assign afi_rdata[62] = hphy_inst_AFIRDATA_bus[62];
assign afi_rdata[63] = hphy_inst_AFIRDATA_bus[63];
assign afi_rdata[64] = hphy_inst_AFIRDATA_bus[64];
assign afi_rdata[65] = hphy_inst_AFIRDATA_bus[65];
assign afi_rdata[66] = hphy_inst_AFIRDATA_bus[66];
assign afi_rdata[67] = hphy_inst_AFIRDATA_bus[67];
assign afi_rdata[68] = hphy_inst_AFIRDATA_bus[68];
assign afi_rdata[69] = hphy_inst_AFIRDATA_bus[69];
assign afi_rdata[70] = hphy_inst_AFIRDATA_bus[70];
assign afi_rdata[71] = hphy_inst_AFIRDATA_bus[71];
assign afi_rdata[72] = hphy_inst_AFIRDATA_bus[72];
assign afi_rdata[73] = hphy_inst_AFIRDATA_bus[73];
assign afi_rdata[74] = hphy_inst_AFIRDATA_bus[74];
assign afi_rdata[75] = hphy_inst_AFIRDATA_bus[75];
assign afi_rdata[76] = hphy_inst_AFIRDATA_bus[76];
assign afi_rdata[77] = hphy_inst_AFIRDATA_bus[77];
assign afi_rdata[78] = hphy_inst_AFIRDATA_bus[78];
assign afi_rdata[79] = hphy_inst_AFIRDATA_bus[79];

assign afi_wlat[0] = hphy_inst_AFIWLAT_bus[0];
assign afi_wlat[1] = hphy_inst_AFIWLAT_bus[1];
assign afi_wlat[2] = hphy_inst_AFIWLAT_bus[2];
assign afi_wlat[3] = hphy_inst_AFIWLAT_bus[3];

assign \phy_ddio_address[0]  = hphy_inst_PHYDDIOADDRDOUT_bus[0];
assign \phy_ddio_address[1]  = hphy_inst_PHYDDIOADDRDOUT_bus[1];
assign \phy_ddio_address[2]  = hphy_inst_PHYDDIOADDRDOUT_bus[2];
assign \phy_ddio_address[3]  = hphy_inst_PHYDDIOADDRDOUT_bus[3];
assign \phy_ddio_address[4]  = hphy_inst_PHYDDIOADDRDOUT_bus[4];
assign \phy_ddio_address[5]  = hphy_inst_PHYDDIOADDRDOUT_bus[5];
assign \phy_ddio_address[6]  = hphy_inst_PHYDDIOADDRDOUT_bus[6];
assign \phy_ddio_address[7]  = hphy_inst_PHYDDIOADDRDOUT_bus[7];
assign \phy_ddio_address[8]  = hphy_inst_PHYDDIOADDRDOUT_bus[8];
assign \phy_ddio_address[9]  = hphy_inst_PHYDDIOADDRDOUT_bus[9];
assign \phy_ddio_address[10]  = hphy_inst_PHYDDIOADDRDOUT_bus[10];
assign \phy_ddio_address[11]  = hphy_inst_PHYDDIOADDRDOUT_bus[11];
assign \phy_ddio_address[12]  = hphy_inst_PHYDDIOADDRDOUT_bus[12];
assign \phy_ddio_address[13]  = hphy_inst_PHYDDIOADDRDOUT_bus[13];
assign \phy_ddio_address[14]  = hphy_inst_PHYDDIOADDRDOUT_bus[14];
assign \phy_ddio_address[15]  = hphy_inst_PHYDDIOADDRDOUT_bus[15];
assign \phy_ddio_address[16]  = hphy_inst_PHYDDIOADDRDOUT_bus[16];
assign \phy_ddio_address[17]  = hphy_inst_PHYDDIOADDRDOUT_bus[17];
assign \phy_ddio_address[18]  = hphy_inst_PHYDDIOADDRDOUT_bus[18];
assign \phy_ddio_address[19]  = hphy_inst_PHYDDIOADDRDOUT_bus[19];
assign \phy_ddio_address[20]  = hphy_inst_PHYDDIOADDRDOUT_bus[20];
assign \phy_ddio_address[21]  = hphy_inst_PHYDDIOADDRDOUT_bus[21];
assign \phy_ddio_address[22]  = hphy_inst_PHYDDIOADDRDOUT_bus[22];
assign \phy_ddio_address[23]  = hphy_inst_PHYDDIOADDRDOUT_bus[23];
assign \phy_ddio_address[24]  = hphy_inst_PHYDDIOADDRDOUT_bus[24];
assign \phy_ddio_address[25]  = hphy_inst_PHYDDIOADDRDOUT_bus[25];
assign \phy_ddio_address[26]  = hphy_inst_PHYDDIOADDRDOUT_bus[26];
assign \phy_ddio_address[27]  = hphy_inst_PHYDDIOADDRDOUT_bus[27];
assign \phy_ddio_address[28]  = hphy_inst_PHYDDIOADDRDOUT_bus[28];
assign \phy_ddio_address[29]  = hphy_inst_PHYDDIOADDRDOUT_bus[29];
assign \phy_ddio_address[30]  = hphy_inst_PHYDDIOADDRDOUT_bus[30];
assign \phy_ddio_address[31]  = hphy_inst_PHYDDIOADDRDOUT_bus[31];
assign \phy_ddio_address[32]  = hphy_inst_PHYDDIOADDRDOUT_bus[32];
assign \phy_ddio_address[33]  = hphy_inst_PHYDDIOADDRDOUT_bus[33];
assign \phy_ddio_address[34]  = hphy_inst_PHYDDIOADDRDOUT_bus[34];
assign \phy_ddio_address[35]  = hphy_inst_PHYDDIOADDRDOUT_bus[35];
assign \phy_ddio_address[36]  = hphy_inst_PHYDDIOADDRDOUT_bus[36];
assign \phy_ddio_address[37]  = hphy_inst_PHYDDIOADDRDOUT_bus[37];
assign \phy_ddio_address[38]  = hphy_inst_PHYDDIOADDRDOUT_bus[38];
assign \phy_ddio_address[39]  = hphy_inst_PHYDDIOADDRDOUT_bus[39];
assign \phy_ddio_address[40]  = hphy_inst_PHYDDIOADDRDOUT_bus[40];
assign \phy_ddio_address[41]  = hphy_inst_PHYDDIOADDRDOUT_bus[41];
assign \phy_ddio_address[42]  = hphy_inst_PHYDDIOADDRDOUT_bus[42];
assign \phy_ddio_address[43]  = hphy_inst_PHYDDIOADDRDOUT_bus[43];
assign \phy_ddio_address[44]  = hphy_inst_PHYDDIOADDRDOUT_bus[44];
assign \phy_ddio_address[45]  = hphy_inst_PHYDDIOADDRDOUT_bus[45];
assign \phy_ddio_address[46]  = hphy_inst_PHYDDIOADDRDOUT_bus[46];
assign \phy_ddio_address[47]  = hphy_inst_PHYDDIOADDRDOUT_bus[47];
assign \phy_ddio_address[48]  = hphy_inst_PHYDDIOADDRDOUT_bus[48];
assign \phy_ddio_address[49]  = hphy_inst_PHYDDIOADDRDOUT_bus[49];
assign \phy_ddio_address[50]  = hphy_inst_PHYDDIOADDRDOUT_bus[50];
assign \phy_ddio_address[51]  = hphy_inst_PHYDDIOADDRDOUT_bus[51];
assign \phy_ddio_address[52]  = hphy_inst_PHYDDIOADDRDOUT_bus[52];
assign \phy_ddio_address[53]  = hphy_inst_PHYDDIOADDRDOUT_bus[53];
assign \phy_ddio_address[54]  = hphy_inst_PHYDDIOADDRDOUT_bus[54];
assign \phy_ddio_address[55]  = hphy_inst_PHYDDIOADDRDOUT_bus[55];
assign \phy_ddio_address[56]  = hphy_inst_PHYDDIOADDRDOUT_bus[56];
assign \phy_ddio_address[57]  = hphy_inst_PHYDDIOADDRDOUT_bus[57];
assign \phy_ddio_address[58]  = hphy_inst_PHYDDIOADDRDOUT_bus[58];
assign \phy_ddio_address[59]  = hphy_inst_PHYDDIOADDRDOUT_bus[59];

assign \phy_ddio_bank[0]  = hphy_inst_PHYDDIOBADOUT_bus[0];
assign \phy_ddio_bank[1]  = hphy_inst_PHYDDIOBADOUT_bus[1];
assign \phy_ddio_bank[2]  = hphy_inst_PHYDDIOBADOUT_bus[2];
assign \phy_ddio_bank[3]  = hphy_inst_PHYDDIOBADOUT_bus[3];
assign \phy_ddio_bank[4]  = hphy_inst_PHYDDIOBADOUT_bus[4];
assign \phy_ddio_bank[5]  = hphy_inst_PHYDDIOBADOUT_bus[5];
assign \phy_ddio_bank[6]  = hphy_inst_PHYDDIOBADOUT_bus[6];
assign \phy_ddio_bank[7]  = hphy_inst_PHYDDIOBADOUT_bus[7];
assign \phy_ddio_bank[8]  = hphy_inst_PHYDDIOBADOUT_bus[8];
assign \phy_ddio_bank[9]  = hphy_inst_PHYDDIOBADOUT_bus[9];
assign \phy_ddio_bank[10]  = hphy_inst_PHYDDIOBADOUT_bus[10];
assign \phy_ddio_bank[11]  = hphy_inst_PHYDDIOBADOUT_bus[11];

assign \phy_ddio_cas_n[0]  = hphy_inst_PHYDDIOCASNDOUT_bus[0];
assign \phy_ddio_cas_n[1]  = hphy_inst_PHYDDIOCASNDOUT_bus[1];
assign \phy_ddio_cas_n[2]  = hphy_inst_PHYDDIOCASNDOUT_bus[2];
assign \phy_ddio_cas_n[3]  = hphy_inst_PHYDDIOCASNDOUT_bus[3];

assign \phy_ddio_ck[0]  = hphy_inst_PHYDDIOCKDOUT_bus[0];
assign \phy_ddio_ck[1]  = hphy_inst_PHYDDIOCKDOUT_bus[1];

assign \phy_ddio_cke[0]  = hphy_inst_PHYDDIOCKEDOUT_bus[0];
assign \phy_ddio_cke[1]  = hphy_inst_PHYDDIOCKEDOUT_bus[1];
assign \phy_ddio_cke[2]  = hphy_inst_PHYDDIOCKEDOUT_bus[2];
assign \phy_ddio_cke[3]  = hphy_inst_PHYDDIOCKEDOUT_bus[3];

assign \phy_ddio_cs_n[0]  = hphy_inst_PHYDDIOCSNDOUT_bus[0];
assign \phy_ddio_cs_n[1]  = hphy_inst_PHYDDIOCSNDOUT_bus[1];
assign \phy_ddio_cs_n[2]  = hphy_inst_PHYDDIOCSNDOUT_bus[2];
assign \phy_ddio_cs_n[3]  = hphy_inst_PHYDDIOCSNDOUT_bus[3];

assign \phy_ddio_dmdout[0]  = hphy_inst_PHYDDIODMDOUT_bus[0];
assign \phy_ddio_dmdout[1]  = hphy_inst_PHYDDIODMDOUT_bus[1];
assign \phy_ddio_dmdout[2]  = hphy_inst_PHYDDIODMDOUT_bus[2];
assign \phy_ddio_dmdout[3]  = hphy_inst_PHYDDIODMDOUT_bus[3];
assign \phy_ddio_dmdout[4]  = hphy_inst_PHYDDIODMDOUT_bus[4];
assign \phy_ddio_dmdout[5]  = hphy_inst_PHYDDIODMDOUT_bus[5];
assign \phy_ddio_dmdout[6]  = hphy_inst_PHYDDIODMDOUT_bus[6];
assign \phy_ddio_dmdout[7]  = hphy_inst_PHYDDIODMDOUT_bus[7];
assign \phy_ddio_dmdout[8]  = hphy_inst_PHYDDIODMDOUT_bus[8];
assign \phy_ddio_dmdout[9]  = hphy_inst_PHYDDIODMDOUT_bus[9];
assign \phy_ddio_dmdout[10]  = hphy_inst_PHYDDIODMDOUT_bus[10];
assign \phy_ddio_dmdout[11]  = hphy_inst_PHYDDIODMDOUT_bus[11];
assign \phy_ddio_dmdout[12]  = hphy_inst_PHYDDIODMDOUT_bus[12];
assign \phy_ddio_dmdout[13]  = hphy_inst_PHYDDIODMDOUT_bus[13];
assign \phy_ddio_dmdout[14]  = hphy_inst_PHYDDIODMDOUT_bus[14];
assign \phy_ddio_dmdout[15]  = hphy_inst_PHYDDIODMDOUT_bus[15];

assign \phy_ddio_dqdout[0]  = hphy_inst_PHYDDIODQDOUT_bus[0];
assign \phy_ddio_dqdout[1]  = hphy_inst_PHYDDIODQDOUT_bus[1];
assign \phy_ddio_dqdout[2]  = hphy_inst_PHYDDIODQDOUT_bus[2];
assign \phy_ddio_dqdout[3]  = hphy_inst_PHYDDIODQDOUT_bus[3];
assign \phy_ddio_dqdout[4]  = hphy_inst_PHYDDIODQDOUT_bus[4];
assign \phy_ddio_dqdout[5]  = hphy_inst_PHYDDIODQDOUT_bus[5];
assign \phy_ddio_dqdout[6]  = hphy_inst_PHYDDIODQDOUT_bus[6];
assign \phy_ddio_dqdout[7]  = hphy_inst_PHYDDIODQDOUT_bus[7];
assign \phy_ddio_dqdout[8]  = hphy_inst_PHYDDIODQDOUT_bus[8];
assign \phy_ddio_dqdout[9]  = hphy_inst_PHYDDIODQDOUT_bus[9];
assign \phy_ddio_dqdout[10]  = hphy_inst_PHYDDIODQDOUT_bus[10];
assign \phy_ddio_dqdout[11]  = hphy_inst_PHYDDIODQDOUT_bus[11];
assign \phy_ddio_dqdout[12]  = hphy_inst_PHYDDIODQDOUT_bus[12];
assign \phy_ddio_dqdout[13]  = hphy_inst_PHYDDIODQDOUT_bus[13];
assign \phy_ddio_dqdout[14]  = hphy_inst_PHYDDIODQDOUT_bus[14];
assign \phy_ddio_dqdout[15]  = hphy_inst_PHYDDIODQDOUT_bus[15];
assign \phy_ddio_dqdout[16]  = hphy_inst_PHYDDIODQDOUT_bus[16];
assign \phy_ddio_dqdout[17]  = hphy_inst_PHYDDIODQDOUT_bus[17];
assign \phy_ddio_dqdout[18]  = hphy_inst_PHYDDIODQDOUT_bus[18];
assign \phy_ddio_dqdout[19]  = hphy_inst_PHYDDIODQDOUT_bus[19];
assign \phy_ddio_dqdout[20]  = hphy_inst_PHYDDIODQDOUT_bus[20];
assign \phy_ddio_dqdout[21]  = hphy_inst_PHYDDIODQDOUT_bus[21];
assign \phy_ddio_dqdout[22]  = hphy_inst_PHYDDIODQDOUT_bus[22];
assign \phy_ddio_dqdout[23]  = hphy_inst_PHYDDIODQDOUT_bus[23];
assign \phy_ddio_dqdout[24]  = hphy_inst_PHYDDIODQDOUT_bus[24];
assign \phy_ddio_dqdout[25]  = hphy_inst_PHYDDIODQDOUT_bus[25];
assign \phy_ddio_dqdout[26]  = hphy_inst_PHYDDIODQDOUT_bus[26];
assign \phy_ddio_dqdout[27]  = hphy_inst_PHYDDIODQDOUT_bus[27];
assign \phy_ddio_dqdout[28]  = hphy_inst_PHYDDIODQDOUT_bus[28];
assign \phy_ddio_dqdout[29]  = hphy_inst_PHYDDIODQDOUT_bus[29];
assign \phy_ddio_dqdout[30]  = hphy_inst_PHYDDIODQDOUT_bus[30];
assign \phy_ddio_dqdout[31]  = hphy_inst_PHYDDIODQDOUT_bus[31];
assign \phy_ddio_dqdout[36]  = hphy_inst_PHYDDIODQDOUT_bus[36];
assign \phy_ddio_dqdout[37]  = hphy_inst_PHYDDIODQDOUT_bus[37];
assign \phy_ddio_dqdout[38]  = hphy_inst_PHYDDIODQDOUT_bus[38];
assign \phy_ddio_dqdout[39]  = hphy_inst_PHYDDIODQDOUT_bus[39];
assign \phy_ddio_dqdout[40]  = hphy_inst_PHYDDIODQDOUT_bus[40];
assign \phy_ddio_dqdout[41]  = hphy_inst_PHYDDIODQDOUT_bus[41];
assign \phy_ddio_dqdout[42]  = hphy_inst_PHYDDIODQDOUT_bus[42];
assign \phy_ddio_dqdout[43]  = hphy_inst_PHYDDIODQDOUT_bus[43];
assign \phy_ddio_dqdout[44]  = hphy_inst_PHYDDIODQDOUT_bus[44];
assign \phy_ddio_dqdout[45]  = hphy_inst_PHYDDIODQDOUT_bus[45];
assign \phy_ddio_dqdout[46]  = hphy_inst_PHYDDIODQDOUT_bus[46];
assign \phy_ddio_dqdout[47]  = hphy_inst_PHYDDIODQDOUT_bus[47];
assign \phy_ddio_dqdout[48]  = hphy_inst_PHYDDIODQDOUT_bus[48];
assign \phy_ddio_dqdout[49]  = hphy_inst_PHYDDIODQDOUT_bus[49];
assign \phy_ddio_dqdout[50]  = hphy_inst_PHYDDIODQDOUT_bus[50];
assign \phy_ddio_dqdout[51]  = hphy_inst_PHYDDIODQDOUT_bus[51];
assign \phy_ddio_dqdout[52]  = hphy_inst_PHYDDIODQDOUT_bus[52];
assign \phy_ddio_dqdout[53]  = hphy_inst_PHYDDIODQDOUT_bus[53];
assign \phy_ddio_dqdout[54]  = hphy_inst_PHYDDIODQDOUT_bus[54];
assign \phy_ddio_dqdout[55]  = hphy_inst_PHYDDIODQDOUT_bus[55];
assign \phy_ddio_dqdout[56]  = hphy_inst_PHYDDIODQDOUT_bus[56];
assign \phy_ddio_dqdout[57]  = hphy_inst_PHYDDIODQDOUT_bus[57];
assign \phy_ddio_dqdout[58]  = hphy_inst_PHYDDIODQDOUT_bus[58];
assign \phy_ddio_dqdout[59]  = hphy_inst_PHYDDIODQDOUT_bus[59];
assign \phy_ddio_dqdout[60]  = hphy_inst_PHYDDIODQDOUT_bus[60];
assign \phy_ddio_dqdout[61]  = hphy_inst_PHYDDIODQDOUT_bus[61];
assign \phy_ddio_dqdout[62]  = hphy_inst_PHYDDIODQDOUT_bus[62];
assign \phy_ddio_dqdout[63]  = hphy_inst_PHYDDIODQDOUT_bus[63];
assign \phy_ddio_dqdout[64]  = hphy_inst_PHYDDIODQDOUT_bus[64];
assign \phy_ddio_dqdout[65]  = hphy_inst_PHYDDIODQDOUT_bus[65];
assign \phy_ddio_dqdout[66]  = hphy_inst_PHYDDIODQDOUT_bus[66];
assign \phy_ddio_dqdout[67]  = hphy_inst_PHYDDIODQDOUT_bus[67];
assign \phy_ddio_dqdout[72]  = hphy_inst_PHYDDIODQDOUT_bus[72];
assign \phy_ddio_dqdout[73]  = hphy_inst_PHYDDIODQDOUT_bus[73];
assign \phy_ddio_dqdout[74]  = hphy_inst_PHYDDIODQDOUT_bus[74];
assign \phy_ddio_dqdout[75]  = hphy_inst_PHYDDIODQDOUT_bus[75];
assign \phy_ddio_dqdout[76]  = hphy_inst_PHYDDIODQDOUT_bus[76];
assign \phy_ddio_dqdout[77]  = hphy_inst_PHYDDIODQDOUT_bus[77];
assign \phy_ddio_dqdout[78]  = hphy_inst_PHYDDIODQDOUT_bus[78];
assign \phy_ddio_dqdout[79]  = hphy_inst_PHYDDIODQDOUT_bus[79];
assign \phy_ddio_dqdout[80]  = hphy_inst_PHYDDIODQDOUT_bus[80];
assign \phy_ddio_dqdout[81]  = hphy_inst_PHYDDIODQDOUT_bus[81];
assign \phy_ddio_dqdout[82]  = hphy_inst_PHYDDIODQDOUT_bus[82];
assign \phy_ddio_dqdout[83]  = hphy_inst_PHYDDIODQDOUT_bus[83];
assign \phy_ddio_dqdout[84]  = hphy_inst_PHYDDIODQDOUT_bus[84];
assign \phy_ddio_dqdout[85]  = hphy_inst_PHYDDIODQDOUT_bus[85];
assign \phy_ddio_dqdout[86]  = hphy_inst_PHYDDIODQDOUT_bus[86];
assign \phy_ddio_dqdout[87]  = hphy_inst_PHYDDIODQDOUT_bus[87];
assign \phy_ddio_dqdout[88]  = hphy_inst_PHYDDIODQDOUT_bus[88];
assign \phy_ddio_dqdout[89]  = hphy_inst_PHYDDIODQDOUT_bus[89];
assign \phy_ddio_dqdout[90]  = hphy_inst_PHYDDIODQDOUT_bus[90];
assign \phy_ddio_dqdout[91]  = hphy_inst_PHYDDIODQDOUT_bus[91];
assign \phy_ddio_dqdout[92]  = hphy_inst_PHYDDIODQDOUT_bus[92];
assign \phy_ddio_dqdout[93]  = hphy_inst_PHYDDIODQDOUT_bus[93];
assign \phy_ddio_dqdout[94]  = hphy_inst_PHYDDIODQDOUT_bus[94];
assign \phy_ddio_dqdout[95]  = hphy_inst_PHYDDIODQDOUT_bus[95];
assign \phy_ddio_dqdout[96]  = hphy_inst_PHYDDIODQDOUT_bus[96];
assign \phy_ddio_dqdout[97]  = hphy_inst_PHYDDIODQDOUT_bus[97];
assign \phy_ddio_dqdout[98]  = hphy_inst_PHYDDIODQDOUT_bus[98];
assign \phy_ddio_dqdout[99]  = hphy_inst_PHYDDIODQDOUT_bus[99];
assign \phy_ddio_dqdout[100]  = hphy_inst_PHYDDIODQDOUT_bus[100];
assign \phy_ddio_dqdout[101]  = hphy_inst_PHYDDIODQDOUT_bus[101];
assign \phy_ddio_dqdout[102]  = hphy_inst_PHYDDIODQDOUT_bus[102];
assign \phy_ddio_dqdout[103]  = hphy_inst_PHYDDIODQDOUT_bus[103];
assign \phy_ddio_dqdout[108]  = hphy_inst_PHYDDIODQDOUT_bus[108];
assign \phy_ddio_dqdout[109]  = hphy_inst_PHYDDIODQDOUT_bus[109];
assign \phy_ddio_dqdout[110]  = hphy_inst_PHYDDIODQDOUT_bus[110];
assign \phy_ddio_dqdout[111]  = hphy_inst_PHYDDIODQDOUT_bus[111];
assign \phy_ddio_dqdout[112]  = hphy_inst_PHYDDIODQDOUT_bus[112];
assign \phy_ddio_dqdout[113]  = hphy_inst_PHYDDIODQDOUT_bus[113];
assign \phy_ddio_dqdout[114]  = hphy_inst_PHYDDIODQDOUT_bus[114];
assign \phy_ddio_dqdout[115]  = hphy_inst_PHYDDIODQDOUT_bus[115];
assign \phy_ddio_dqdout[116]  = hphy_inst_PHYDDIODQDOUT_bus[116];
assign \phy_ddio_dqdout[117]  = hphy_inst_PHYDDIODQDOUT_bus[117];
assign \phy_ddio_dqdout[118]  = hphy_inst_PHYDDIODQDOUT_bus[118];
assign \phy_ddio_dqdout[119]  = hphy_inst_PHYDDIODQDOUT_bus[119];
assign \phy_ddio_dqdout[120]  = hphy_inst_PHYDDIODQDOUT_bus[120];
assign \phy_ddio_dqdout[121]  = hphy_inst_PHYDDIODQDOUT_bus[121];
assign \phy_ddio_dqdout[122]  = hphy_inst_PHYDDIODQDOUT_bus[122];
assign \phy_ddio_dqdout[123]  = hphy_inst_PHYDDIODQDOUT_bus[123];
assign \phy_ddio_dqdout[124]  = hphy_inst_PHYDDIODQDOUT_bus[124];
assign \phy_ddio_dqdout[125]  = hphy_inst_PHYDDIODQDOUT_bus[125];
assign \phy_ddio_dqdout[126]  = hphy_inst_PHYDDIODQDOUT_bus[126];
assign \phy_ddio_dqdout[127]  = hphy_inst_PHYDDIODQDOUT_bus[127];
assign \phy_ddio_dqdout[128]  = hphy_inst_PHYDDIODQDOUT_bus[128];
assign \phy_ddio_dqdout[129]  = hphy_inst_PHYDDIODQDOUT_bus[129];
assign \phy_ddio_dqdout[130]  = hphy_inst_PHYDDIODQDOUT_bus[130];
assign \phy_ddio_dqdout[131]  = hphy_inst_PHYDDIODQDOUT_bus[131];
assign \phy_ddio_dqdout[132]  = hphy_inst_PHYDDIODQDOUT_bus[132];
assign \phy_ddio_dqdout[133]  = hphy_inst_PHYDDIODQDOUT_bus[133];
assign \phy_ddio_dqdout[134]  = hphy_inst_PHYDDIODQDOUT_bus[134];
assign \phy_ddio_dqdout[135]  = hphy_inst_PHYDDIODQDOUT_bus[135];
assign \phy_ddio_dqdout[136]  = hphy_inst_PHYDDIODQDOUT_bus[136];
assign \phy_ddio_dqdout[137]  = hphy_inst_PHYDDIODQDOUT_bus[137];
assign \phy_ddio_dqdout[138]  = hphy_inst_PHYDDIODQDOUT_bus[138];
assign \phy_ddio_dqdout[139]  = hphy_inst_PHYDDIODQDOUT_bus[139];

assign \phy_ddio_dqoe[0]  = hphy_inst_PHYDDIODQOE_bus[0];
assign \phy_ddio_dqoe[1]  = hphy_inst_PHYDDIODQOE_bus[1];
assign \phy_ddio_dqoe[2]  = hphy_inst_PHYDDIODQOE_bus[2];
assign \phy_ddio_dqoe[3]  = hphy_inst_PHYDDIODQOE_bus[3];
assign \phy_ddio_dqoe[4]  = hphy_inst_PHYDDIODQOE_bus[4];
assign \phy_ddio_dqoe[5]  = hphy_inst_PHYDDIODQOE_bus[5];
assign \phy_ddio_dqoe[6]  = hphy_inst_PHYDDIODQOE_bus[6];
assign \phy_ddio_dqoe[7]  = hphy_inst_PHYDDIODQOE_bus[7];
assign \phy_ddio_dqoe[8]  = hphy_inst_PHYDDIODQOE_bus[8];
assign \phy_ddio_dqoe[9]  = hphy_inst_PHYDDIODQOE_bus[9];
assign \phy_ddio_dqoe[10]  = hphy_inst_PHYDDIODQOE_bus[10];
assign \phy_ddio_dqoe[11]  = hphy_inst_PHYDDIODQOE_bus[11];
assign \phy_ddio_dqoe[12]  = hphy_inst_PHYDDIODQOE_bus[12];
assign \phy_ddio_dqoe[13]  = hphy_inst_PHYDDIODQOE_bus[13];
assign \phy_ddio_dqoe[14]  = hphy_inst_PHYDDIODQOE_bus[14];
assign \phy_ddio_dqoe[15]  = hphy_inst_PHYDDIODQOE_bus[15];
assign \phy_ddio_dqoe[18]  = hphy_inst_PHYDDIODQOE_bus[18];
assign \phy_ddio_dqoe[19]  = hphy_inst_PHYDDIODQOE_bus[19];
assign \phy_ddio_dqoe[20]  = hphy_inst_PHYDDIODQOE_bus[20];
assign \phy_ddio_dqoe[21]  = hphy_inst_PHYDDIODQOE_bus[21];
assign \phy_ddio_dqoe[22]  = hphy_inst_PHYDDIODQOE_bus[22];
assign \phy_ddio_dqoe[23]  = hphy_inst_PHYDDIODQOE_bus[23];
assign \phy_ddio_dqoe[24]  = hphy_inst_PHYDDIODQOE_bus[24];
assign \phy_ddio_dqoe[25]  = hphy_inst_PHYDDIODQOE_bus[25];
assign \phy_ddio_dqoe[26]  = hphy_inst_PHYDDIODQOE_bus[26];
assign \phy_ddio_dqoe[27]  = hphy_inst_PHYDDIODQOE_bus[27];
assign \phy_ddio_dqoe[28]  = hphy_inst_PHYDDIODQOE_bus[28];
assign \phy_ddio_dqoe[29]  = hphy_inst_PHYDDIODQOE_bus[29];
assign \phy_ddio_dqoe[30]  = hphy_inst_PHYDDIODQOE_bus[30];
assign \phy_ddio_dqoe[31]  = hphy_inst_PHYDDIODQOE_bus[31];
assign \phy_ddio_dqoe[32]  = hphy_inst_PHYDDIODQOE_bus[32];
assign \phy_ddio_dqoe[33]  = hphy_inst_PHYDDIODQOE_bus[33];
assign \phy_ddio_dqoe[36]  = hphy_inst_PHYDDIODQOE_bus[36];
assign \phy_ddio_dqoe[37]  = hphy_inst_PHYDDIODQOE_bus[37];
assign \phy_ddio_dqoe[38]  = hphy_inst_PHYDDIODQOE_bus[38];
assign \phy_ddio_dqoe[39]  = hphy_inst_PHYDDIODQOE_bus[39];
assign \phy_ddio_dqoe[40]  = hphy_inst_PHYDDIODQOE_bus[40];
assign \phy_ddio_dqoe[41]  = hphy_inst_PHYDDIODQOE_bus[41];
assign \phy_ddio_dqoe[42]  = hphy_inst_PHYDDIODQOE_bus[42];
assign \phy_ddio_dqoe[43]  = hphy_inst_PHYDDIODQOE_bus[43];
assign \phy_ddio_dqoe[44]  = hphy_inst_PHYDDIODQOE_bus[44];
assign \phy_ddio_dqoe[45]  = hphy_inst_PHYDDIODQOE_bus[45];
assign \phy_ddio_dqoe[46]  = hphy_inst_PHYDDIODQOE_bus[46];
assign \phy_ddio_dqoe[47]  = hphy_inst_PHYDDIODQOE_bus[47];
assign \phy_ddio_dqoe[48]  = hphy_inst_PHYDDIODQOE_bus[48];
assign \phy_ddio_dqoe[49]  = hphy_inst_PHYDDIODQOE_bus[49];
assign \phy_ddio_dqoe[50]  = hphy_inst_PHYDDIODQOE_bus[50];
assign \phy_ddio_dqoe[51]  = hphy_inst_PHYDDIODQOE_bus[51];
assign \phy_ddio_dqoe[54]  = hphy_inst_PHYDDIODQOE_bus[54];
assign \phy_ddio_dqoe[55]  = hphy_inst_PHYDDIODQOE_bus[55];
assign \phy_ddio_dqoe[56]  = hphy_inst_PHYDDIODQOE_bus[56];
assign \phy_ddio_dqoe[57]  = hphy_inst_PHYDDIODQOE_bus[57];
assign \phy_ddio_dqoe[58]  = hphy_inst_PHYDDIODQOE_bus[58];
assign \phy_ddio_dqoe[59]  = hphy_inst_PHYDDIODQOE_bus[59];
assign \phy_ddio_dqoe[60]  = hphy_inst_PHYDDIODQOE_bus[60];
assign \phy_ddio_dqoe[61]  = hphy_inst_PHYDDIODQOE_bus[61];
assign \phy_ddio_dqoe[62]  = hphy_inst_PHYDDIODQOE_bus[62];
assign \phy_ddio_dqoe[63]  = hphy_inst_PHYDDIODQOE_bus[63];
assign \phy_ddio_dqoe[64]  = hphy_inst_PHYDDIODQOE_bus[64];
assign \phy_ddio_dqoe[65]  = hphy_inst_PHYDDIODQOE_bus[65];
assign \phy_ddio_dqoe[66]  = hphy_inst_PHYDDIODQOE_bus[66];
assign \phy_ddio_dqoe[67]  = hphy_inst_PHYDDIODQOE_bus[67];
assign \phy_ddio_dqoe[68]  = hphy_inst_PHYDDIODQOE_bus[68];
assign \phy_ddio_dqoe[69]  = hphy_inst_PHYDDIODQOE_bus[69];

assign \phy_ddio_dqs_dout[0]  = hphy_inst_PHYDDIODQSDOUT_bus[0];
assign \phy_ddio_dqs_dout[1]  = hphy_inst_PHYDDIODQSDOUT_bus[1];
assign \phy_ddio_dqs_dout[2]  = hphy_inst_PHYDDIODQSDOUT_bus[2];
assign \phy_ddio_dqs_dout[3]  = hphy_inst_PHYDDIODQSDOUT_bus[3];
assign \phy_ddio_dqs_dout[4]  = hphy_inst_PHYDDIODQSDOUT_bus[4];
assign \phy_ddio_dqs_dout[5]  = hphy_inst_PHYDDIODQSDOUT_bus[5];
assign \phy_ddio_dqs_dout[6]  = hphy_inst_PHYDDIODQSDOUT_bus[6];
assign \phy_ddio_dqs_dout[7]  = hphy_inst_PHYDDIODQSDOUT_bus[7];
assign \phy_ddio_dqs_dout[8]  = hphy_inst_PHYDDIODQSDOUT_bus[8];
assign \phy_ddio_dqs_dout[9]  = hphy_inst_PHYDDIODQSDOUT_bus[9];
assign \phy_ddio_dqs_dout[10]  = hphy_inst_PHYDDIODQSDOUT_bus[10];
assign \phy_ddio_dqs_dout[11]  = hphy_inst_PHYDDIODQSDOUT_bus[11];
assign \phy_ddio_dqs_dout[12]  = hphy_inst_PHYDDIODQSDOUT_bus[12];
assign \phy_ddio_dqs_dout[13]  = hphy_inst_PHYDDIODQSDOUT_bus[13];
assign \phy_ddio_dqs_dout[14]  = hphy_inst_PHYDDIODQSDOUT_bus[14];
assign \phy_ddio_dqs_dout[15]  = hphy_inst_PHYDDIODQSDOUT_bus[15];

assign \phy_ddio_dqslogic_aclr_fifoctrl[0]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[0];
assign \phy_ddio_dqslogic_aclr_fifoctrl[1]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[1];
assign \phy_ddio_dqslogic_aclr_fifoctrl[2]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[2];
assign \phy_ddio_dqslogic_aclr_fifoctrl[3]  = hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus[3];

assign \phy_ddio_dqslogic_aclr_pstamble[0]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[0];
assign \phy_ddio_dqslogic_aclr_pstamble[1]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[1];
assign \phy_ddio_dqslogic_aclr_pstamble[2]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[2];
assign \phy_ddio_dqslogic_aclr_pstamble[3]  = hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus[3];

assign \phy_ddio_dqslogic_dqsena[0]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[0];
assign \phy_ddio_dqslogic_dqsena[1]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[1];
assign \phy_ddio_dqslogic_dqsena[2]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[2];
assign \phy_ddio_dqslogic_dqsena[3]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[3];
assign \phy_ddio_dqslogic_dqsena[4]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[4];
assign \phy_ddio_dqslogic_dqsena[5]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[5];
assign \phy_ddio_dqslogic_dqsena[6]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[6];
assign \phy_ddio_dqslogic_dqsena[7]  = hphy_inst_PHYDDIODQSLOGICDQSENA_bus[7];

assign \phy_ddio_dqslogic_fiforeset[0]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[0];
assign \phy_ddio_dqslogic_fiforeset[1]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[1];
assign \phy_ddio_dqslogic_fiforeset[2]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[2];
assign \phy_ddio_dqslogic_fiforeset[3]  = hphy_inst_PHYDDIODQSLOGICFIFORESET_bus[3];

assign \phy_ddio_dqslogic_incrdataen[0]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[0];
assign \phy_ddio_dqslogic_incrdataen[1]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[1];
assign \phy_ddio_dqslogic_incrdataen[2]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[2];
assign \phy_ddio_dqslogic_incrdataen[3]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[3];
assign \phy_ddio_dqslogic_incrdataen[4]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[4];
assign \phy_ddio_dqslogic_incrdataen[5]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[5];
assign \phy_ddio_dqslogic_incrdataen[6]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[6];
assign \phy_ddio_dqslogic_incrdataen[7]  = hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus[7];

assign \phy_ddio_dqslogic_incwrptr[0]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[0];
assign \phy_ddio_dqslogic_incwrptr[1]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[1];
assign \phy_ddio_dqslogic_incwrptr[2]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[2];
assign \phy_ddio_dqslogic_incwrptr[3]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[3];
assign \phy_ddio_dqslogic_incwrptr[4]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[4];
assign \phy_ddio_dqslogic_incwrptr[5]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[5];
assign \phy_ddio_dqslogic_incwrptr[6]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[6];
assign \phy_ddio_dqslogic_incwrptr[7]  = hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus[7];

assign \phy_ddio_dqslogic_oct[0]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[0];
assign \phy_ddio_dqslogic_oct[1]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[1];
assign \phy_ddio_dqslogic_oct[2]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[2];
assign \phy_ddio_dqslogic_oct[3]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[3];
assign \phy_ddio_dqslogic_oct[4]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[4];
assign \phy_ddio_dqslogic_oct[5]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[5];
assign \phy_ddio_dqslogic_oct[6]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[6];
assign \phy_ddio_dqslogic_oct[7]  = hphy_inst_PHYDDIODQSLOGICOCT_bus[7];

assign \phy_ddio_dqslogic_readlatency[0]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[0];
assign \phy_ddio_dqslogic_readlatency[1]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[1];
assign \phy_ddio_dqslogic_readlatency[2]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[2];
assign \phy_ddio_dqslogic_readlatency[3]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[3];
assign \phy_ddio_dqslogic_readlatency[4]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[4];
assign \phy_ddio_dqslogic_readlatency[5]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[5];
assign \phy_ddio_dqslogic_readlatency[6]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[6];
assign \phy_ddio_dqslogic_readlatency[7]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[7];
assign \phy_ddio_dqslogic_readlatency[8]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[8];
assign \phy_ddio_dqslogic_readlatency[9]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[9];
assign \phy_ddio_dqslogic_readlatency[10]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[10];
assign \phy_ddio_dqslogic_readlatency[11]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[11];
assign \phy_ddio_dqslogic_readlatency[12]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[12];
assign \phy_ddio_dqslogic_readlatency[13]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[13];
assign \phy_ddio_dqslogic_readlatency[14]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[14];
assign \phy_ddio_dqslogic_readlatency[15]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[15];
assign \phy_ddio_dqslogic_readlatency[16]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[16];
assign \phy_ddio_dqslogic_readlatency[17]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[17];
assign \phy_ddio_dqslogic_readlatency[18]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[18];
assign \phy_ddio_dqslogic_readlatency[19]  = hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus[19];

assign \phy_ddio_dqs_oe[0]  = hphy_inst_PHYDDIODQSOE_bus[0];
assign \phy_ddio_dqs_oe[1]  = hphy_inst_PHYDDIODQSOE_bus[1];
assign \phy_ddio_dqs_oe[2]  = hphy_inst_PHYDDIODQSOE_bus[2];
assign \phy_ddio_dqs_oe[3]  = hphy_inst_PHYDDIODQSOE_bus[3];
assign \phy_ddio_dqs_oe[4]  = hphy_inst_PHYDDIODQSOE_bus[4];
assign \phy_ddio_dqs_oe[5]  = hphy_inst_PHYDDIODQSOE_bus[5];
assign \phy_ddio_dqs_oe[6]  = hphy_inst_PHYDDIODQSOE_bus[6];
assign \phy_ddio_dqs_oe[7]  = hphy_inst_PHYDDIODQSOE_bus[7];

assign \phy_ddio_odt[0]  = hphy_inst_PHYDDIOODTDOUT_bus[0];
assign \phy_ddio_odt[1]  = hphy_inst_PHYDDIOODTDOUT_bus[1];
assign \phy_ddio_odt[2]  = hphy_inst_PHYDDIOODTDOUT_bus[2];
assign \phy_ddio_odt[3]  = hphy_inst_PHYDDIOODTDOUT_bus[3];

assign \phy_ddio_ras_n[0]  = hphy_inst_PHYDDIORASNDOUT_bus[0];
assign \phy_ddio_ras_n[1]  = hphy_inst_PHYDDIORASNDOUT_bus[1];
assign \phy_ddio_ras_n[2]  = hphy_inst_PHYDDIORASNDOUT_bus[2];
assign \phy_ddio_ras_n[3]  = hphy_inst_PHYDDIORASNDOUT_bus[3];

assign \phy_ddio_reset_n[0]  = hphy_inst_PHYDDIORESETNDOUT_bus[0];
assign \phy_ddio_reset_n[1]  = hphy_inst_PHYDDIORESETNDOUT_bus[1];
assign \phy_ddio_reset_n[2]  = hphy_inst_PHYDDIORESETNDOUT_bus[2];
assign \phy_ddio_reset_n[3]  = hphy_inst_PHYDDIORESETNDOUT_bus[3];

assign \phy_ddio_we_n[0]  = hphy_inst_PHYDDIOWENDOUT_bus[0];
assign \phy_ddio_we_n[1]  = hphy_inst_PHYDDIOWENDOUT_bus[1];
assign \phy_ddio_we_n[2]  = hphy_inst_PHYDDIOWENDOUT_bus[2];
assign \phy_ddio_we_n[3]  = hphy_inst_PHYDDIOWENDOUT_bus[3];

terminal_qsys_hps_sdram_p0_acv_hard_io_pads uio_pads(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.dqsin1(dqsin1),
	.pad_gen0raw_input1(pad_gen0raw_input1),
	.pad_gen1raw_input1(pad_gen1raw_input1),
	.pad_gen2raw_input1(pad_gen2raw_input1),
	.pad_gen3raw_input1(pad_gen3raw_input1),
	.pad_gen4raw_input1(pad_gen4raw_input1),
	.pad_gen5raw_input1(pad_gen5raw_input1),
	.pad_gen6raw_input1(pad_gen6raw_input1),
	.pad_gen7raw_input1(pad_gen7raw_input1),
	.dqsin2(dqsin2),
	.pad_gen0raw_input2(pad_gen0raw_input2),
	.pad_gen1raw_input2(pad_gen1raw_input2),
	.pad_gen2raw_input2(pad_gen2raw_input2),
	.pad_gen3raw_input2(pad_gen3raw_input2),
	.pad_gen4raw_input2(pad_gen4raw_input2),
	.pad_gen5raw_input2(pad_gen5raw_input2),
	.pad_gen6raw_input2(pad_gen6raw_input2),
	.pad_gen7raw_input2(pad_gen7raw_input2),
	.dqsin3(dqsin3),
	.pad_gen0raw_input3(pad_gen0raw_input3),
	.pad_gen1raw_input3(pad_gen1raw_input3),
	.pad_gen2raw_input3(pad_gen2raw_input3),
	.pad_gen3raw_input3(pad_gen3raw_input3),
	.pad_gen4raw_input3(pad_gen4raw_input3),
	.pad_gen5raw_input3(pad_gen5raw_input3),
	.pad_gen6raw_input3(pad_gen6raw_input3),
	.pad_gen7raw_input3(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_output_pad_gen0delayed_data_out1(extra_output_pad_gen0delayed_data_out1),
	.extra_output_pad_gen0delayed_data_out2(extra_output_pad_gen0delayed_data_out2),
	.extra_output_pad_gen0delayed_data_out3(extra_output_pad_gen0delayed_data_out3),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(\phy_ddio_address[0] ),
	.phy_ddio_address_1(\phy_ddio_address[1] ),
	.phy_ddio_address_2(\phy_ddio_address[2] ),
	.phy_ddio_address_3(\phy_ddio_address[3] ),
	.phy_ddio_address_4(\phy_ddio_address[4] ),
	.phy_ddio_address_5(\phy_ddio_address[5] ),
	.phy_ddio_address_6(\phy_ddio_address[6] ),
	.phy_ddio_address_7(\phy_ddio_address[7] ),
	.phy_ddio_address_8(\phy_ddio_address[8] ),
	.phy_ddio_address_9(\phy_ddio_address[9] ),
	.phy_ddio_address_10(\phy_ddio_address[10] ),
	.phy_ddio_address_11(\phy_ddio_address[11] ),
	.phy_ddio_address_12(\phy_ddio_address[12] ),
	.phy_ddio_address_13(\phy_ddio_address[13] ),
	.phy_ddio_address_14(\phy_ddio_address[14] ),
	.phy_ddio_address_15(\phy_ddio_address[15] ),
	.phy_ddio_address_16(\phy_ddio_address[16] ),
	.phy_ddio_address_17(\phy_ddio_address[17] ),
	.phy_ddio_address_18(\phy_ddio_address[18] ),
	.phy_ddio_address_19(\phy_ddio_address[19] ),
	.phy_ddio_address_20(\phy_ddio_address[20] ),
	.phy_ddio_address_21(\phy_ddio_address[21] ),
	.phy_ddio_address_22(\phy_ddio_address[22] ),
	.phy_ddio_address_23(\phy_ddio_address[23] ),
	.phy_ddio_address_24(\phy_ddio_address[24] ),
	.phy_ddio_address_25(\phy_ddio_address[25] ),
	.phy_ddio_address_26(\phy_ddio_address[26] ),
	.phy_ddio_address_27(\phy_ddio_address[27] ),
	.phy_ddio_address_28(\phy_ddio_address[28] ),
	.phy_ddio_address_29(\phy_ddio_address[29] ),
	.phy_ddio_address_30(\phy_ddio_address[30] ),
	.phy_ddio_address_31(\phy_ddio_address[31] ),
	.phy_ddio_address_32(\phy_ddio_address[32] ),
	.phy_ddio_address_33(\phy_ddio_address[33] ),
	.phy_ddio_address_34(\phy_ddio_address[34] ),
	.phy_ddio_address_35(\phy_ddio_address[35] ),
	.phy_ddio_address_36(\phy_ddio_address[36] ),
	.phy_ddio_address_37(\phy_ddio_address[37] ),
	.phy_ddio_address_38(\phy_ddio_address[38] ),
	.phy_ddio_address_39(\phy_ddio_address[39] ),
	.phy_ddio_address_40(\phy_ddio_address[40] ),
	.phy_ddio_address_41(\phy_ddio_address[41] ),
	.phy_ddio_address_42(\phy_ddio_address[42] ),
	.phy_ddio_address_43(\phy_ddio_address[43] ),
	.phy_ddio_address_44(\phy_ddio_address[44] ),
	.phy_ddio_address_45(\phy_ddio_address[45] ),
	.phy_ddio_address_46(\phy_ddio_address[46] ),
	.phy_ddio_address_47(\phy_ddio_address[47] ),
	.phy_ddio_address_48(\phy_ddio_address[48] ),
	.phy_ddio_address_49(\phy_ddio_address[49] ),
	.phy_ddio_address_50(\phy_ddio_address[50] ),
	.phy_ddio_address_51(\phy_ddio_address[51] ),
	.phy_ddio_address_52(\phy_ddio_address[52] ),
	.phy_ddio_address_53(\phy_ddio_address[53] ),
	.phy_ddio_address_54(\phy_ddio_address[54] ),
	.phy_ddio_address_55(\phy_ddio_address[55] ),
	.phy_ddio_address_56(\phy_ddio_address[56] ),
	.phy_ddio_address_57(\phy_ddio_address[57] ),
	.phy_ddio_address_58(\phy_ddio_address[58] ),
	.phy_ddio_address_59(\phy_ddio_address[59] ),
	.phy_ddio_bank_0(\phy_ddio_bank[0] ),
	.phy_ddio_bank_1(\phy_ddio_bank[1] ),
	.phy_ddio_bank_2(\phy_ddio_bank[2] ),
	.phy_ddio_bank_3(\phy_ddio_bank[3] ),
	.phy_ddio_bank_4(\phy_ddio_bank[4] ),
	.phy_ddio_bank_5(\phy_ddio_bank[5] ),
	.phy_ddio_bank_6(\phy_ddio_bank[6] ),
	.phy_ddio_bank_7(\phy_ddio_bank[7] ),
	.phy_ddio_bank_8(\phy_ddio_bank[8] ),
	.phy_ddio_bank_9(\phy_ddio_bank[9] ),
	.phy_ddio_bank_10(\phy_ddio_bank[10] ),
	.phy_ddio_bank_11(\phy_ddio_bank[11] ),
	.phy_ddio_cas_n_0(\phy_ddio_cas_n[0] ),
	.phy_ddio_cas_n_1(\phy_ddio_cas_n[1] ),
	.phy_ddio_cas_n_2(\phy_ddio_cas_n[2] ),
	.phy_ddio_cas_n_3(\phy_ddio_cas_n[3] ),
	.phy_ddio_ck_0(\phy_ddio_ck[0] ),
	.phy_ddio_ck_1(\phy_ddio_ck[1] ),
	.phy_ddio_cke_0(\phy_ddio_cke[0] ),
	.phy_ddio_cke_1(\phy_ddio_cke[1] ),
	.phy_ddio_cke_2(\phy_ddio_cke[2] ),
	.phy_ddio_cke_3(\phy_ddio_cke[3] ),
	.phy_ddio_cs_n_0(\phy_ddio_cs_n[0] ),
	.phy_ddio_cs_n_1(\phy_ddio_cs_n[1] ),
	.phy_ddio_cs_n_2(\phy_ddio_cs_n[2] ),
	.phy_ddio_cs_n_3(\phy_ddio_cs_n[3] ),
	.phy_ddio_dmdout_0(\phy_ddio_dmdout[0] ),
	.phy_ddio_dmdout_1(\phy_ddio_dmdout[1] ),
	.phy_ddio_dmdout_2(\phy_ddio_dmdout[2] ),
	.phy_ddio_dmdout_3(\phy_ddio_dmdout[3] ),
	.phy_ddio_dmdout_4(\phy_ddio_dmdout[4] ),
	.phy_ddio_dmdout_5(\phy_ddio_dmdout[5] ),
	.phy_ddio_dmdout_6(\phy_ddio_dmdout[6] ),
	.phy_ddio_dmdout_7(\phy_ddio_dmdout[7] ),
	.phy_ddio_dmdout_8(\phy_ddio_dmdout[8] ),
	.phy_ddio_dmdout_9(\phy_ddio_dmdout[9] ),
	.phy_ddio_dmdout_10(\phy_ddio_dmdout[10] ),
	.phy_ddio_dmdout_11(\phy_ddio_dmdout[11] ),
	.phy_ddio_dmdout_12(\phy_ddio_dmdout[12] ),
	.phy_ddio_dmdout_13(\phy_ddio_dmdout[13] ),
	.phy_ddio_dmdout_14(\phy_ddio_dmdout[14] ),
	.phy_ddio_dmdout_15(\phy_ddio_dmdout[15] ),
	.phy_ddio_dqdout_0(\phy_ddio_dqdout[0] ),
	.phy_ddio_dqdout_1(\phy_ddio_dqdout[1] ),
	.phy_ddio_dqdout_2(\phy_ddio_dqdout[2] ),
	.phy_ddio_dqdout_3(\phy_ddio_dqdout[3] ),
	.phy_ddio_dqdout_4(\phy_ddio_dqdout[4] ),
	.phy_ddio_dqdout_5(\phy_ddio_dqdout[5] ),
	.phy_ddio_dqdout_6(\phy_ddio_dqdout[6] ),
	.phy_ddio_dqdout_7(\phy_ddio_dqdout[7] ),
	.phy_ddio_dqdout_8(\phy_ddio_dqdout[8] ),
	.phy_ddio_dqdout_9(\phy_ddio_dqdout[9] ),
	.phy_ddio_dqdout_10(\phy_ddio_dqdout[10] ),
	.phy_ddio_dqdout_11(\phy_ddio_dqdout[11] ),
	.phy_ddio_dqdout_12(\phy_ddio_dqdout[12] ),
	.phy_ddio_dqdout_13(\phy_ddio_dqdout[13] ),
	.phy_ddio_dqdout_14(\phy_ddio_dqdout[14] ),
	.phy_ddio_dqdout_15(\phy_ddio_dqdout[15] ),
	.phy_ddio_dqdout_16(\phy_ddio_dqdout[16] ),
	.phy_ddio_dqdout_17(\phy_ddio_dqdout[17] ),
	.phy_ddio_dqdout_18(\phy_ddio_dqdout[18] ),
	.phy_ddio_dqdout_19(\phy_ddio_dqdout[19] ),
	.phy_ddio_dqdout_20(\phy_ddio_dqdout[20] ),
	.phy_ddio_dqdout_21(\phy_ddio_dqdout[21] ),
	.phy_ddio_dqdout_22(\phy_ddio_dqdout[22] ),
	.phy_ddio_dqdout_23(\phy_ddio_dqdout[23] ),
	.phy_ddio_dqdout_24(\phy_ddio_dqdout[24] ),
	.phy_ddio_dqdout_25(\phy_ddio_dqdout[25] ),
	.phy_ddio_dqdout_26(\phy_ddio_dqdout[26] ),
	.phy_ddio_dqdout_27(\phy_ddio_dqdout[27] ),
	.phy_ddio_dqdout_28(\phy_ddio_dqdout[28] ),
	.phy_ddio_dqdout_29(\phy_ddio_dqdout[29] ),
	.phy_ddio_dqdout_30(\phy_ddio_dqdout[30] ),
	.phy_ddio_dqdout_31(\phy_ddio_dqdout[31] ),
	.phy_ddio_dqdout_36(\phy_ddio_dqdout[36] ),
	.phy_ddio_dqdout_37(\phy_ddio_dqdout[37] ),
	.phy_ddio_dqdout_38(\phy_ddio_dqdout[38] ),
	.phy_ddio_dqdout_39(\phy_ddio_dqdout[39] ),
	.phy_ddio_dqdout_40(\phy_ddio_dqdout[40] ),
	.phy_ddio_dqdout_41(\phy_ddio_dqdout[41] ),
	.phy_ddio_dqdout_42(\phy_ddio_dqdout[42] ),
	.phy_ddio_dqdout_43(\phy_ddio_dqdout[43] ),
	.phy_ddio_dqdout_44(\phy_ddio_dqdout[44] ),
	.phy_ddio_dqdout_45(\phy_ddio_dqdout[45] ),
	.phy_ddio_dqdout_46(\phy_ddio_dqdout[46] ),
	.phy_ddio_dqdout_47(\phy_ddio_dqdout[47] ),
	.phy_ddio_dqdout_48(\phy_ddio_dqdout[48] ),
	.phy_ddio_dqdout_49(\phy_ddio_dqdout[49] ),
	.phy_ddio_dqdout_50(\phy_ddio_dqdout[50] ),
	.phy_ddio_dqdout_51(\phy_ddio_dqdout[51] ),
	.phy_ddio_dqdout_52(\phy_ddio_dqdout[52] ),
	.phy_ddio_dqdout_53(\phy_ddio_dqdout[53] ),
	.phy_ddio_dqdout_54(\phy_ddio_dqdout[54] ),
	.phy_ddio_dqdout_55(\phy_ddio_dqdout[55] ),
	.phy_ddio_dqdout_56(\phy_ddio_dqdout[56] ),
	.phy_ddio_dqdout_57(\phy_ddio_dqdout[57] ),
	.phy_ddio_dqdout_58(\phy_ddio_dqdout[58] ),
	.phy_ddio_dqdout_59(\phy_ddio_dqdout[59] ),
	.phy_ddio_dqdout_60(\phy_ddio_dqdout[60] ),
	.phy_ddio_dqdout_61(\phy_ddio_dqdout[61] ),
	.phy_ddio_dqdout_62(\phy_ddio_dqdout[62] ),
	.phy_ddio_dqdout_63(\phy_ddio_dqdout[63] ),
	.phy_ddio_dqdout_64(\phy_ddio_dqdout[64] ),
	.phy_ddio_dqdout_65(\phy_ddio_dqdout[65] ),
	.phy_ddio_dqdout_66(\phy_ddio_dqdout[66] ),
	.phy_ddio_dqdout_67(\phy_ddio_dqdout[67] ),
	.phy_ddio_dqdout_72(\phy_ddio_dqdout[72] ),
	.phy_ddio_dqdout_73(\phy_ddio_dqdout[73] ),
	.phy_ddio_dqdout_74(\phy_ddio_dqdout[74] ),
	.phy_ddio_dqdout_75(\phy_ddio_dqdout[75] ),
	.phy_ddio_dqdout_76(\phy_ddio_dqdout[76] ),
	.phy_ddio_dqdout_77(\phy_ddio_dqdout[77] ),
	.phy_ddio_dqdout_78(\phy_ddio_dqdout[78] ),
	.phy_ddio_dqdout_79(\phy_ddio_dqdout[79] ),
	.phy_ddio_dqdout_80(\phy_ddio_dqdout[80] ),
	.phy_ddio_dqdout_81(\phy_ddio_dqdout[81] ),
	.phy_ddio_dqdout_82(\phy_ddio_dqdout[82] ),
	.phy_ddio_dqdout_83(\phy_ddio_dqdout[83] ),
	.phy_ddio_dqdout_84(\phy_ddio_dqdout[84] ),
	.phy_ddio_dqdout_85(\phy_ddio_dqdout[85] ),
	.phy_ddio_dqdout_86(\phy_ddio_dqdout[86] ),
	.phy_ddio_dqdout_87(\phy_ddio_dqdout[87] ),
	.phy_ddio_dqdout_88(\phy_ddio_dqdout[88] ),
	.phy_ddio_dqdout_89(\phy_ddio_dqdout[89] ),
	.phy_ddio_dqdout_90(\phy_ddio_dqdout[90] ),
	.phy_ddio_dqdout_91(\phy_ddio_dqdout[91] ),
	.phy_ddio_dqdout_92(\phy_ddio_dqdout[92] ),
	.phy_ddio_dqdout_93(\phy_ddio_dqdout[93] ),
	.phy_ddio_dqdout_94(\phy_ddio_dqdout[94] ),
	.phy_ddio_dqdout_95(\phy_ddio_dqdout[95] ),
	.phy_ddio_dqdout_96(\phy_ddio_dqdout[96] ),
	.phy_ddio_dqdout_97(\phy_ddio_dqdout[97] ),
	.phy_ddio_dqdout_98(\phy_ddio_dqdout[98] ),
	.phy_ddio_dqdout_99(\phy_ddio_dqdout[99] ),
	.phy_ddio_dqdout_100(\phy_ddio_dqdout[100] ),
	.phy_ddio_dqdout_101(\phy_ddio_dqdout[101] ),
	.phy_ddio_dqdout_102(\phy_ddio_dqdout[102] ),
	.phy_ddio_dqdout_103(\phy_ddio_dqdout[103] ),
	.phy_ddio_dqdout_108(\phy_ddio_dqdout[108] ),
	.phy_ddio_dqdout_109(\phy_ddio_dqdout[109] ),
	.phy_ddio_dqdout_110(\phy_ddio_dqdout[110] ),
	.phy_ddio_dqdout_111(\phy_ddio_dqdout[111] ),
	.phy_ddio_dqdout_112(\phy_ddio_dqdout[112] ),
	.phy_ddio_dqdout_113(\phy_ddio_dqdout[113] ),
	.phy_ddio_dqdout_114(\phy_ddio_dqdout[114] ),
	.phy_ddio_dqdout_115(\phy_ddio_dqdout[115] ),
	.phy_ddio_dqdout_116(\phy_ddio_dqdout[116] ),
	.phy_ddio_dqdout_117(\phy_ddio_dqdout[117] ),
	.phy_ddio_dqdout_118(\phy_ddio_dqdout[118] ),
	.phy_ddio_dqdout_119(\phy_ddio_dqdout[119] ),
	.phy_ddio_dqdout_120(\phy_ddio_dqdout[120] ),
	.phy_ddio_dqdout_121(\phy_ddio_dqdout[121] ),
	.phy_ddio_dqdout_122(\phy_ddio_dqdout[122] ),
	.phy_ddio_dqdout_123(\phy_ddio_dqdout[123] ),
	.phy_ddio_dqdout_124(\phy_ddio_dqdout[124] ),
	.phy_ddio_dqdout_125(\phy_ddio_dqdout[125] ),
	.phy_ddio_dqdout_126(\phy_ddio_dqdout[126] ),
	.phy_ddio_dqdout_127(\phy_ddio_dqdout[127] ),
	.phy_ddio_dqdout_128(\phy_ddio_dqdout[128] ),
	.phy_ddio_dqdout_129(\phy_ddio_dqdout[129] ),
	.phy_ddio_dqdout_130(\phy_ddio_dqdout[130] ),
	.phy_ddio_dqdout_131(\phy_ddio_dqdout[131] ),
	.phy_ddio_dqdout_132(\phy_ddio_dqdout[132] ),
	.phy_ddio_dqdout_133(\phy_ddio_dqdout[133] ),
	.phy_ddio_dqdout_134(\phy_ddio_dqdout[134] ),
	.phy_ddio_dqdout_135(\phy_ddio_dqdout[135] ),
	.phy_ddio_dqdout_136(\phy_ddio_dqdout[136] ),
	.phy_ddio_dqdout_137(\phy_ddio_dqdout[137] ),
	.phy_ddio_dqdout_138(\phy_ddio_dqdout[138] ),
	.phy_ddio_dqdout_139(\phy_ddio_dqdout[139] ),
	.phy_ddio_dqoe_0(\phy_ddio_dqoe[0] ),
	.phy_ddio_dqoe_1(\phy_ddio_dqoe[1] ),
	.phy_ddio_dqoe_2(\phy_ddio_dqoe[2] ),
	.phy_ddio_dqoe_3(\phy_ddio_dqoe[3] ),
	.phy_ddio_dqoe_4(\phy_ddio_dqoe[4] ),
	.phy_ddio_dqoe_5(\phy_ddio_dqoe[5] ),
	.phy_ddio_dqoe_6(\phy_ddio_dqoe[6] ),
	.phy_ddio_dqoe_7(\phy_ddio_dqoe[7] ),
	.phy_ddio_dqoe_8(\phy_ddio_dqoe[8] ),
	.phy_ddio_dqoe_9(\phy_ddio_dqoe[9] ),
	.phy_ddio_dqoe_10(\phy_ddio_dqoe[10] ),
	.phy_ddio_dqoe_11(\phy_ddio_dqoe[11] ),
	.phy_ddio_dqoe_12(\phy_ddio_dqoe[12] ),
	.phy_ddio_dqoe_13(\phy_ddio_dqoe[13] ),
	.phy_ddio_dqoe_14(\phy_ddio_dqoe[14] ),
	.phy_ddio_dqoe_15(\phy_ddio_dqoe[15] ),
	.phy_ddio_dqoe_18(\phy_ddio_dqoe[18] ),
	.phy_ddio_dqoe_19(\phy_ddio_dqoe[19] ),
	.phy_ddio_dqoe_20(\phy_ddio_dqoe[20] ),
	.phy_ddio_dqoe_21(\phy_ddio_dqoe[21] ),
	.phy_ddio_dqoe_22(\phy_ddio_dqoe[22] ),
	.phy_ddio_dqoe_23(\phy_ddio_dqoe[23] ),
	.phy_ddio_dqoe_24(\phy_ddio_dqoe[24] ),
	.phy_ddio_dqoe_25(\phy_ddio_dqoe[25] ),
	.phy_ddio_dqoe_26(\phy_ddio_dqoe[26] ),
	.phy_ddio_dqoe_27(\phy_ddio_dqoe[27] ),
	.phy_ddio_dqoe_28(\phy_ddio_dqoe[28] ),
	.phy_ddio_dqoe_29(\phy_ddio_dqoe[29] ),
	.phy_ddio_dqoe_30(\phy_ddio_dqoe[30] ),
	.phy_ddio_dqoe_31(\phy_ddio_dqoe[31] ),
	.phy_ddio_dqoe_32(\phy_ddio_dqoe[32] ),
	.phy_ddio_dqoe_33(\phy_ddio_dqoe[33] ),
	.phy_ddio_dqoe_36(\phy_ddio_dqoe[36] ),
	.phy_ddio_dqoe_37(\phy_ddio_dqoe[37] ),
	.phy_ddio_dqoe_38(\phy_ddio_dqoe[38] ),
	.phy_ddio_dqoe_39(\phy_ddio_dqoe[39] ),
	.phy_ddio_dqoe_40(\phy_ddio_dqoe[40] ),
	.phy_ddio_dqoe_41(\phy_ddio_dqoe[41] ),
	.phy_ddio_dqoe_42(\phy_ddio_dqoe[42] ),
	.phy_ddio_dqoe_43(\phy_ddio_dqoe[43] ),
	.phy_ddio_dqoe_44(\phy_ddio_dqoe[44] ),
	.phy_ddio_dqoe_45(\phy_ddio_dqoe[45] ),
	.phy_ddio_dqoe_46(\phy_ddio_dqoe[46] ),
	.phy_ddio_dqoe_47(\phy_ddio_dqoe[47] ),
	.phy_ddio_dqoe_48(\phy_ddio_dqoe[48] ),
	.phy_ddio_dqoe_49(\phy_ddio_dqoe[49] ),
	.phy_ddio_dqoe_50(\phy_ddio_dqoe[50] ),
	.phy_ddio_dqoe_51(\phy_ddio_dqoe[51] ),
	.phy_ddio_dqoe_54(\phy_ddio_dqoe[54] ),
	.phy_ddio_dqoe_55(\phy_ddio_dqoe[55] ),
	.phy_ddio_dqoe_56(\phy_ddio_dqoe[56] ),
	.phy_ddio_dqoe_57(\phy_ddio_dqoe[57] ),
	.phy_ddio_dqoe_58(\phy_ddio_dqoe[58] ),
	.phy_ddio_dqoe_59(\phy_ddio_dqoe[59] ),
	.phy_ddio_dqoe_60(\phy_ddio_dqoe[60] ),
	.phy_ddio_dqoe_61(\phy_ddio_dqoe[61] ),
	.phy_ddio_dqoe_62(\phy_ddio_dqoe[62] ),
	.phy_ddio_dqoe_63(\phy_ddio_dqoe[63] ),
	.phy_ddio_dqoe_64(\phy_ddio_dqoe[64] ),
	.phy_ddio_dqoe_65(\phy_ddio_dqoe[65] ),
	.phy_ddio_dqoe_66(\phy_ddio_dqoe[66] ),
	.phy_ddio_dqoe_67(\phy_ddio_dqoe[67] ),
	.phy_ddio_dqoe_68(\phy_ddio_dqoe[68] ),
	.phy_ddio_dqoe_69(\phy_ddio_dqoe[69] ),
	.phy_ddio_dqs_dout_0(\phy_ddio_dqs_dout[0] ),
	.phy_ddio_dqs_dout_1(\phy_ddio_dqs_dout[1] ),
	.phy_ddio_dqs_dout_2(\phy_ddio_dqs_dout[2] ),
	.phy_ddio_dqs_dout_3(\phy_ddio_dqs_dout[3] ),
	.phy_ddio_dqs_dout_4(\phy_ddio_dqs_dout[4] ),
	.phy_ddio_dqs_dout_5(\phy_ddio_dqs_dout[5] ),
	.phy_ddio_dqs_dout_6(\phy_ddio_dqs_dout[6] ),
	.phy_ddio_dqs_dout_7(\phy_ddio_dqs_dout[7] ),
	.phy_ddio_dqs_dout_8(\phy_ddio_dqs_dout[8] ),
	.phy_ddio_dqs_dout_9(\phy_ddio_dqs_dout[9] ),
	.phy_ddio_dqs_dout_10(\phy_ddio_dqs_dout[10] ),
	.phy_ddio_dqs_dout_11(\phy_ddio_dqs_dout[11] ),
	.phy_ddio_dqs_dout_12(\phy_ddio_dqs_dout[12] ),
	.phy_ddio_dqs_dout_13(\phy_ddio_dqs_dout[13] ),
	.phy_ddio_dqs_dout_14(\phy_ddio_dqs_dout[14] ),
	.phy_ddio_dqs_dout_15(\phy_ddio_dqs_dout[15] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(\phy_ddio_dqslogic_aclr_fifoctrl[0] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(\phy_ddio_dqslogic_aclr_fifoctrl[1] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(\phy_ddio_dqslogic_aclr_fifoctrl[2] ),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(\phy_ddio_dqslogic_aclr_fifoctrl[3] ),
	.phy_ddio_dqslogic_aclr_pstamble_0(\phy_ddio_dqslogic_aclr_pstamble[0] ),
	.phy_ddio_dqslogic_aclr_pstamble_1(\phy_ddio_dqslogic_aclr_pstamble[1] ),
	.phy_ddio_dqslogic_aclr_pstamble_2(\phy_ddio_dqslogic_aclr_pstamble[2] ),
	.phy_ddio_dqslogic_aclr_pstamble_3(\phy_ddio_dqslogic_aclr_pstamble[3] ),
	.phy_ddio_dqslogic_dqsena_0(\phy_ddio_dqslogic_dqsena[0] ),
	.phy_ddio_dqslogic_dqsena_1(\phy_ddio_dqslogic_dqsena[1] ),
	.phy_ddio_dqslogic_dqsena_2(\phy_ddio_dqslogic_dqsena[2] ),
	.phy_ddio_dqslogic_dqsena_3(\phy_ddio_dqslogic_dqsena[3] ),
	.phy_ddio_dqslogic_dqsena_4(\phy_ddio_dqslogic_dqsena[4] ),
	.phy_ddio_dqslogic_dqsena_5(\phy_ddio_dqslogic_dqsena[5] ),
	.phy_ddio_dqslogic_dqsena_6(\phy_ddio_dqslogic_dqsena[6] ),
	.phy_ddio_dqslogic_dqsena_7(\phy_ddio_dqslogic_dqsena[7] ),
	.phy_ddio_dqslogic_fiforeset_0(\phy_ddio_dqslogic_fiforeset[0] ),
	.phy_ddio_dqslogic_fiforeset_1(\phy_ddio_dqslogic_fiforeset[1] ),
	.phy_ddio_dqslogic_fiforeset_2(\phy_ddio_dqslogic_fiforeset[2] ),
	.phy_ddio_dqslogic_fiforeset_3(\phy_ddio_dqslogic_fiforeset[3] ),
	.phy_ddio_dqslogic_incrdataen_0(\phy_ddio_dqslogic_incrdataen[0] ),
	.phy_ddio_dqslogic_incrdataen_1(\phy_ddio_dqslogic_incrdataen[1] ),
	.phy_ddio_dqslogic_incrdataen_2(\phy_ddio_dqslogic_incrdataen[2] ),
	.phy_ddio_dqslogic_incrdataen_3(\phy_ddio_dqslogic_incrdataen[3] ),
	.phy_ddio_dqslogic_incrdataen_4(\phy_ddio_dqslogic_incrdataen[4] ),
	.phy_ddio_dqslogic_incrdataen_5(\phy_ddio_dqslogic_incrdataen[5] ),
	.phy_ddio_dqslogic_incrdataen_6(\phy_ddio_dqslogic_incrdataen[6] ),
	.phy_ddio_dqslogic_incrdataen_7(\phy_ddio_dqslogic_incrdataen[7] ),
	.phy_ddio_dqslogic_incwrptr_0(\phy_ddio_dqslogic_incwrptr[0] ),
	.phy_ddio_dqslogic_incwrptr_1(\phy_ddio_dqslogic_incwrptr[1] ),
	.phy_ddio_dqslogic_incwrptr_2(\phy_ddio_dqslogic_incwrptr[2] ),
	.phy_ddio_dqslogic_incwrptr_3(\phy_ddio_dqslogic_incwrptr[3] ),
	.phy_ddio_dqslogic_incwrptr_4(\phy_ddio_dqslogic_incwrptr[4] ),
	.phy_ddio_dqslogic_incwrptr_5(\phy_ddio_dqslogic_incwrptr[5] ),
	.phy_ddio_dqslogic_incwrptr_6(\phy_ddio_dqslogic_incwrptr[6] ),
	.phy_ddio_dqslogic_incwrptr_7(\phy_ddio_dqslogic_incwrptr[7] ),
	.phy_ddio_dqslogic_oct_0(\phy_ddio_dqslogic_oct[0] ),
	.phy_ddio_dqslogic_oct_1(\phy_ddio_dqslogic_oct[1] ),
	.phy_ddio_dqslogic_oct_2(\phy_ddio_dqslogic_oct[2] ),
	.phy_ddio_dqslogic_oct_3(\phy_ddio_dqslogic_oct[3] ),
	.phy_ddio_dqslogic_oct_4(\phy_ddio_dqslogic_oct[4] ),
	.phy_ddio_dqslogic_oct_5(\phy_ddio_dqslogic_oct[5] ),
	.phy_ddio_dqslogic_oct_6(\phy_ddio_dqslogic_oct[6] ),
	.phy_ddio_dqslogic_oct_7(\phy_ddio_dqslogic_oct[7] ),
	.phy_ddio_dqslogic_readlatency_0(\phy_ddio_dqslogic_readlatency[0] ),
	.phy_ddio_dqslogic_readlatency_1(\phy_ddio_dqslogic_readlatency[1] ),
	.phy_ddio_dqslogic_readlatency_2(\phy_ddio_dqslogic_readlatency[2] ),
	.phy_ddio_dqslogic_readlatency_3(\phy_ddio_dqslogic_readlatency[3] ),
	.phy_ddio_dqslogic_readlatency_4(\phy_ddio_dqslogic_readlatency[4] ),
	.phy_ddio_dqslogic_readlatency_5(\phy_ddio_dqslogic_readlatency[5] ),
	.phy_ddio_dqslogic_readlatency_6(\phy_ddio_dqslogic_readlatency[6] ),
	.phy_ddio_dqslogic_readlatency_7(\phy_ddio_dqslogic_readlatency[7] ),
	.phy_ddio_dqslogic_readlatency_8(\phy_ddio_dqslogic_readlatency[8] ),
	.phy_ddio_dqslogic_readlatency_9(\phy_ddio_dqslogic_readlatency[9] ),
	.phy_ddio_dqslogic_readlatency_10(\phy_ddio_dqslogic_readlatency[10] ),
	.phy_ddio_dqslogic_readlatency_11(\phy_ddio_dqslogic_readlatency[11] ),
	.phy_ddio_dqslogic_readlatency_12(\phy_ddio_dqslogic_readlatency[12] ),
	.phy_ddio_dqslogic_readlatency_13(\phy_ddio_dqslogic_readlatency[13] ),
	.phy_ddio_dqslogic_readlatency_14(\phy_ddio_dqslogic_readlatency[14] ),
	.phy_ddio_dqslogic_readlatency_15(\phy_ddio_dqslogic_readlatency[15] ),
	.phy_ddio_dqslogic_readlatency_16(\phy_ddio_dqslogic_readlatency[16] ),
	.phy_ddio_dqslogic_readlatency_17(\phy_ddio_dqslogic_readlatency[17] ),
	.phy_ddio_dqslogic_readlatency_18(\phy_ddio_dqslogic_readlatency[18] ),
	.phy_ddio_dqslogic_readlatency_19(\phy_ddio_dqslogic_readlatency[19] ),
	.phy_ddio_dqs_oe_0(\phy_ddio_dqs_oe[0] ),
	.phy_ddio_dqs_oe_1(\phy_ddio_dqs_oe[1] ),
	.phy_ddio_dqs_oe_2(\phy_ddio_dqs_oe[2] ),
	.phy_ddio_dqs_oe_3(\phy_ddio_dqs_oe[3] ),
	.phy_ddio_dqs_oe_4(\phy_ddio_dqs_oe[4] ),
	.phy_ddio_dqs_oe_5(\phy_ddio_dqs_oe[5] ),
	.phy_ddio_dqs_oe_6(\phy_ddio_dqs_oe[6] ),
	.phy_ddio_dqs_oe_7(\phy_ddio_dqs_oe[7] ),
	.phy_ddio_odt_0(\phy_ddio_odt[0] ),
	.phy_ddio_odt_1(\phy_ddio_odt[1] ),
	.phy_ddio_odt_2(\phy_ddio_odt[2] ),
	.phy_ddio_odt_3(\phy_ddio_odt[3] ),
	.phy_ddio_ras_n_0(\phy_ddio_ras_n[0] ),
	.phy_ddio_ras_n_1(\phy_ddio_ras_n[1] ),
	.phy_ddio_ras_n_2(\phy_ddio_ras_n[2] ),
	.phy_ddio_ras_n_3(\phy_ddio_ras_n[3] ),
	.phy_ddio_reset_n_0(\phy_ddio_reset_n[0] ),
	.phy_ddio_reset_n_1(\phy_ddio_reset_n[1] ),
	.phy_ddio_reset_n_2(\phy_ddio_reset_n[2] ),
	.phy_ddio_reset_n_3(\phy_ddio_reset_n[3] ),
	.phy_ddio_we_n_0(\phy_ddio_we_n[0] ),
	.phy_ddio_we_n_1(\phy_ddio_we_n[1] ),
	.phy_ddio_we_n_2(\phy_ddio_we_n[2] ),
	.phy_ddio_we_n_3(\phy_ddio_we_n[3] ),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.pad_gen0delayed_data_out1(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_11(pad_gen0delayed_oe_11),
	.delayed_oct1(delayed_oct1),
	.pad_gen1delayed_data_out1(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_11(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out1(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_11(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out1(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_11(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out1(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_11(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out1(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_11(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out1(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_11(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out1(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_11(pad_gen7delayed_oe_11),
	.pad_gen0delayed_data_out2(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_12(pad_gen0delayed_oe_12),
	.delayed_oct2(delayed_oct2),
	.pad_gen1delayed_data_out2(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_12(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out2(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_12(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out2(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_12(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out2(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_12(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out2(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_12(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out2(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_12(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out2(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_12(pad_gen7delayed_oe_12),
	.pad_gen0delayed_data_out3(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_13(pad_gen0delayed_oe_13),
	.delayed_oct3(delayed_oct3),
	.pad_gen1delayed_data_out3(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_13(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out3(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_13(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out3(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_13(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out3(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_13(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out3(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_13(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out3(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_13(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out3(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_13(pad_gen7delayed_oe_13),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.os1(os1),
	.os_bar1(os_bar1),
	.diff_oe1(diff_oe1),
	.diff_oe_bar1(diff_oe_bar1),
	.diff_dtc1(diff_dtc1),
	.diff_dtc_bar1(diff_dtc_bar1),
	.os2(os2),
	.os_bar2(os_bar2),
	.diff_oe2(diff_oe2),
	.diff_oe_bar2(diff_oe_bar2),
	.diff_dtc2(diff_dtc2),
	.diff_dtc_bar2(diff_dtc_bar2),
	.os3(os3),
	.os_bar3(os_bar3),
	.diff_oe3(diff_oe3),
	.diff_oe_bar3(diff_oe_bar3),
	.diff_dtc3(diff_dtc3),
	.diff_dtc_bar3(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_0(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_1(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_2(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_3(\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_01(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_11(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_21(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_31(\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_02(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_12(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_22(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_32(\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.input_path_gen0read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ),
	.input_path_gen0read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ),
	.input_path_gen0read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ),
	.input_path_gen0read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ),
	.input_path_gen1read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ),
	.input_path_gen1read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ),
	.input_path_gen1read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ),
	.input_path_gen1read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ),
	.input_path_gen2read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ),
	.input_path_gen2read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ),
	.input_path_gen2read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ),
	.input_path_gen2read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ),
	.input_path_gen3read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ),
	.input_path_gen3read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ),
	.input_path_gen3read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ),
	.input_path_gen3read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ),
	.input_path_gen4read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ),
	.input_path_gen4read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ),
	.input_path_gen4read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ),
	.input_path_gen4read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ),
	.input_path_gen5read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ),
	.input_path_gen5read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ),
	.input_path_gen5read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ),
	.input_path_gen5read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ),
	.input_path_gen6read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ),
	.input_path_gen6read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ),
	.input_path_gen6read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ),
	.input_path_gen6read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ),
	.input_path_gen7read_fifo_out_03(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ),
	.input_path_gen7read_fifo_out_13(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ),
	.input_path_gen7read_fifo_out_23(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ),
	.input_path_gen7read_fifo_out_33(\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ),
	.ddio_phy_dqslogic_rdatavalid({ddio_phy_dqslogic_rdatavalid_unconnected_wire_4,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

terminal_qsys_hps_sdram_p0_acv_ldc_25 memphy_ldc(
	.pll_dqs_clk(afi_clk),
	.pll_hr_clk(afi_clk),
	.afi_clk(ctl_clk),
	.avl_clk(\memphy_ldc|leveled_hr_clocks[0] ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_mem_phy hphy_inst(
	.aficasn(afi_cas_n[0]),
	.afimemclkdisable(afi_mem_clk_disable[0]),
	.afirasn(afi_ras_n[0]),
	.afirstn(afi_rst_n[0]),
	.afiwen(afi_we_n[0]),
	.avlread(gnd),
	.avlresetn(gnd),
	.avlwrite(gnd),
	.globalresetn(gnd),
	.iointcasnaclr(gnd),
	.iointrasnaclr(gnd),
	.iointresetnaclr(gnd),
	.iointwenaclr(gnd),
	.plladdrcmdclk(!ctl_clk),
	.pllaficlk(ctl_clk),
	.pllavlclk(\memphy_ldc|leveled_hr_clocks[0] ),
	.plllocked(gnd),
	.scanen(gnd),
	.softresetn(gnd),
	.afiaddr({afi_addr[19],afi_addr[18],afi_addr[17],afi_addr[16],afi_addr[15],afi_addr[14],afi_addr[13],afi_addr[12],afi_addr[11],afi_addr[10],afi_addr[9],afi_addr[8],afi_addr[7],afi_addr[6],afi_addr[5],afi_addr[4],afi_addr[3],afi_addr[2],afi_addr[1],afi_addr[0]}),
	.afiba({afi_ba[2],afi_ba[1],afi_ba[0]}),
	.aficke({afi_cke[1],afi_cke[0]}),
	.aficsn({afi_cs_n[1],afi_cs_n[0]}),
	.afidm({afi_dm[9],afi_dm[8],afi_dm[7],afi_dm[6],afi_dm[5],afi_dm[4],afi_dm[3],afi_dm[2],afi_dm[1],afi_dm[0]}),
	.afidqsburst({afi_dqs_burst[4],afi_dqs_burst[3],afi_dqs_burst[2],afi_dqs_burst[1],afi_dqs_burst[0]}),
	.afiodt({afi_odt[1],afi_odt[0]}),
	.afirdataen({afi_rdata_en[4],afi_rdata_en[3],afi_rdata_en[2],afi_rdata_en[1],afi_rdata_en[0]}),
	.afirdataenfull({afi_rdata_en_full[4],afi_rdata_en_full[3],afi_rdata_en_full[2],afi_rdata_en_full[1],afi_rdata_en_full[0]}),
	.afiwdata({afi_wdata[79],afi_wdata[78],afi_wdata[77],afi_wdata[76],afi_wdata[75],afi_wdata[74],afi_wdata[73],afi_wdata[72],afi_wdata[71],afi_wdata[70],afi_wdata[69],afi_wdata[68],afi_wdata[67],afi_wdata[66],afi_wdata[65],afi_wdata[64],afi_wdata[63],afi_wdata[62],afi_wdata[61],afi_wdata[60],afi_wdata[59],afi_wdata[58],afi_wdata[57],afi_wdata[56],afi_wdata[55],afi_wdata[54],afi_wdata[53],afi_wdata[52],
afi_wdata[51],afi_wdata[50],afi_wdata[49],afi_wdata[48],afi_wdata[47],afi_wdata[46],afi_wdata[45],afi_wdata[44],afi_wdata[43],afi_wdata[42],afi_wdata[41],afi_wdata[40],afi_wdata[39],afi_wdata[38],afi_wdata[37],afi_wdata[36],afi_wdata[35],afi_wdata[34],afi_wdata[33],afi_wdata[32],afi_wdata[31],afi_wdata[30],afi_wdata[29],afi_wdata[28],afi_wdata[27],afi_wdata[26],afi_wdata[25],afi_wdata[24],
afi_wdata[23],afi_wdata[22],afi_wdata[21],afi_wdata[20],afi_wdata[19],afi_wdata[18],afi_wdata[17],afi_wdata[16],afi_wdata[15],afi_wdata[14],afi_wdata[13],afi_wdata[12],afi_wdata[11],afi_wdata[10],afi_wdata[9],afi_wdata[8],afi_wdata[7],afi_wdata[6],afi_wdata[5],afi_wdata[4],afi_wdata[3],afi_wdata[2],afi_wdata[1],afi_wdata[0]}),
	.afiwdatavalid({afi_wdata_valid[4],afi_wdata_valid[3],afi_wdata_valid[2],afi_wdata_valid[1],afi_wdata_valid[0]}),
	.avladdress({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.avlwritedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cfgaddlat({gnd,gnd,gnd,cfg_addlat[4],cfg_addlat[3],cfg_addlat[2],cfg_addlat[1],cfg_addlat[0]}),
	.cfgbankaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_bankaddrwidth[2],cfg_bankaddrwidth[1],cfg_bankaddrwidth[0]}),
	.cfgcaswrlat({gnd,gnd,gnd,gnd,cfg_caswrlat[3],cfg_caswrlat[2],cfg_caswrlat[1],cfg_caswrlat[0]}),
	.cfgcoladdrwidth({gnd,gnd,gnd,cfg_coladdrwidth[4],cfg_coladdrwidth[3],cfg_coladdrwidth[2],cfg_coladdrwidth[1],cfg_coladdrwidth[0]}),
	.cfgcsaddrwidth({gnd,gnd,gnd,gnd,gnd,cfg_csaddrwidth[2],cfg_csaddrwidth[1],cfg_csaddrwidth[0]}),
	.cfgdevicewidth({gnd,gnd,gnd,gnd,cfg_devicewidth[3],cfg_devicewidth[2],cfg_devicewidth[1],cfg_devicewidth[0]}),
	.cfgdramconfig({gnd,gnd,gnd,cfg_dramconfig[20],cfg_dramconfig[19],cfg_dramconfig[18],cfg_dramconfig[17],cfg_dramconfig[16],cfg_dramconfig[15],cfg_dramconfig[14],cfg_dramconfig[13],cfg_dramconfig[12],cfg_dramconfig[11],cfg_dramconfig[10],cfg_dramconfig[9],cfg_dramconfig[8],cfg_dramconfig[7],cfg_dramconfig[6],cfg_dramconfig[5],cfg_dramconfig[4],
cfg_dramconfig[3],cfg_dramconfig[2],cfg_dramconfig[1],cfg_dramconfig[0]}),
	.cfginterfacewidth({cfg_interfacewidth[7],cfg_interfacewidth[6],cfg_interfacewidth[5],cfg_interfacewidth[4],cfg_interfacewidth[3],cfg_interfacewidth[2],cfg_interfacewidth[1],cfg_interfacewidth[0]}),
	.cfgrowaddrwidth({gnd,gnd,gnd,cfg_rowaddrwidth[4],cfg_rowaddrwidth[3],cfg_rowaddrwidth[2],cfg_rowaddrwidth[1],cfg_rowaddrwidth[0]}),
	.cfgtcl({gnd,gnd,gnd,cfg_tcl[4],cfg_tcl[3],cfg_tcl[2],cfg_tcl[1],cfg_tcl[0]}),
	.cfgtmrd({gnd,gnd,gnd,gnd,cfg_tmrd[3],cfg_tmrd[2],cfg_tmrd[1],cfg_tmrd[0]}),
	.cfgtrefi({gnd,gnd,gnd,cfg_trefi[12],cfg_trefi[11],cfg_trefi[10],cfg_trefi[9],cfg_trefi[8],cfg_trefi[7],cfg_trefi[6],cfg_trefi[5],cfg_trefi[4],cfg_trefi[3],cfg_trefi[2],cfg_trefi[1],cfg_trefi[0]}),
	.cfgtrfc({cfg_trfc[7],cfg_trfc[6],cfg_trfc[5],cfg_trfc[4],cfg_trfc[3],cfg_trfc[2],cfg_trfc[1],cfg_trfc[0]}),
	.cfgtwr({gnd,gnd,gnd,gnd,cfg_twr[3],cfg_twr[2],cfg_twr[1],cfg_twr[0]}),
	.ddiophydqdin({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] ,gnd,gnd,gnd,gnd,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[7].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[6].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[5].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[4].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[3].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[2].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[1].read_fifo_out[0] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[3] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[2] ,\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[1] ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|input_path_gen[0].read_fifo_out[0] }),
	.ddiophydqslogicrdatavalid({vcc,\uio_pads|dq_ddio[3].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[2].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,\uio_pads|dq_ddio[1].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid ,
\uio_pads|dq_ddio[0].ubidir_dq_dqs|altdq_dqs2_inst|lfifo_rdata_valid }),
	.iointaddraclr(16'b0000000000000000),
	.iointaddrdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointbaaclr(3'b000),
	.iointbadout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointcasndout({gnd,gnd,gnd,gnd}),
	.iointckdout({gnd,gnd,gnd,gnd}),
	.iointckeaclr(2'b00),
	.iointckedout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointckndout({gnd,gnd,gnd,gnd}),
	.iointcsnaclr(2'b00),
	.iointcsndout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdmdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd}),
	.iointdqsbdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsboe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicaclrfifoctrl(5'b00000),
	.iointdqslogicaclrpstamble(5'b00000),
	.iointdqslogicdqsena({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicfiforeset({gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincrdataen({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicincwrptr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicoct({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqslogicreadlatency({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointdqsoe({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointodtaclr(2'b00),
	.iointodtdout({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.iointrasndout({gnd,gnd,gnd,gnd}),
	.iointresetndout({gnd,gnd,gnd,gnd}),
	.iointwendout({gnd,gnd,gnd,gnd}),
	.aficalfail(afi_cal_fail),
	.aficalsuccess(afi_cal_success),
	.afirdatavalid(afi_rdata_valid[0]),
	.avlwaitrequest(),
	.ctlresetn(ctl_reset_n),
	.iointaficalfail(),
	.iointaficalsuccess(),
	.phyddiocasnaclr(),
	.phyddiorasnaclr(),
	.phyddioresetnaclr(),
	.phyddiowenaclr(),
	.phyresetn(),
	.afirdata(hphy_inst_AFIRDATA_bus),
	.afirlat(),
	.afiwlat(hphy_inst_AFIWLAT_bus),
	.avlreaddata(),
	.iointafirlat(),
	.iointafiwlat(),
	.iointdqdin(),
	.iointdqslogicrdatavalid(),
	.phyddioaddraclr(),
	.phyddioaddrdout(hphy_inst_PHYDDIOADDRDOUT_bus),
	.phyddiobaaclr(),
	.phyddiobadout(hphy_inst_PHYDDIOBADOUT_bus),
	.phyddiocasndout(hphy_inst_PHYDDIOCASNDOUT_bus),
	.phyddiockdout(hphy_inst_PHYDDIOCKDOUT_bus),
	.phyddiockeaclr(),
	.phyddiockedout(hphy_inst_PHYDDIOCKEDOUT_bus),
	.phyddiockndout(),
	.phyddiocsnaclr(),
	.phyddiocsndout(hphy_inst_PHYDDIOCSNDOUT_bus),
	.phyddiodmdout(hphy_inst_PHYDDIODMDOUT_bus),
	.phyddiodqdout(hphy_inst_PHYDDIODQDOUT_bus),
	.phyddiodqoe(hphy_inst_PHYDDIODQOE_bus),
	.phyddiodqsbdout(),
	.phyddiodqsboe(),
	.phyddiodqsdout(hphy_inst_PHYDDIODQSDOUT_bus),
	.phyddiodqslogicaclrfifoctrl(hphy_inst_PHYDDIODQSLOGICACLRFIFOCTRL_bus),
	.phyddiodqslogicaclrpstamble(hphy_inst_PHYDDIODQSLOGICACLRPSTAMBLE_bus),
	.phyddiodqslogicdqsena(hphy_inst_PHYDDIODQSLOGICDQSENA_bus),
	.phyddiodqslogicfiforeset(hphy_inst_PHYDDIODQSLOGICFIFORESET_bus),
	.phyddiodqslogicincrdataen(hphy_inst_PHYDDIODQSLOGICINCRDATAEN_bus),
	.phyddiodqslogicincwrptr(hphy_inst_PHYDDIODQSLOGICINCWRPTR_bus),
	.phyddiodqslogicoct(hphy_inst_PHYDDIODQSLOGICOCT_bus),
	.phyddiodqslogicreadlatency(hphy_inst_PHYDDIODQSLOGICREADLATENCY_bus),
	.phyddiodqsoe(hphy_inst_PHYDDIODQSOE_bus),
	.phyddioodtaclr(),
	.phyddioodtdout(hphy_inst_PHYDDIOODTDOUT_bus),
	.phyddiorasndout(hphy_inst_PHYDDIORASNDOUT_bus),
	.phyddioresetndout(hphy_inst_PHYDDIORESETNDOUT_bus),
	.phyddiowendout(hphy_inst_PHYDDIOWENDOUT_bus));
defparam hphy_inst.hphy_ac_ddr_disable = "true";
defparam hphy_inst.hphy_atpg_en = "false";
defparam hphy_inst.hphy_csr_pipelineglobalenable = "true";
defparam hphy_inst.hphy_datapath_ac_delay = "one_and_half_cycles";
defparam hphy_inst.hphy_datapath_delay = "one_cycle";
defparam hphy_inst.hphy_reset_delay_en = "false";
defparam hphy_inst.hphy_use_hphy = "true";
defparam hphy_inst.hphy_wrap_back_en = "false";
defparam hphy_inst.m_hphy_ac_rom_content = 1200'b100000011100000000000000000000100000011110000000000000000000010000000010000000010000110001010000000010000000010100110000010000000010010000000001000100010000000010100000000000010000010000000010110000000000000000010000001110000000010000000000010000000010000000010001001001010000000010000000010011001000010000000010100000000000100100010000000010010000000000001000010000000010110000000000000000110000011110000000000000000000111000011110000000000000000000110000011110000000000000000000010000011010000000000000000000010000011010110000000000000000010000001010000000010000000000010000010010000000000000000000011100100110000000000000000000011100100110110000000000000000011100100110000000000000001000011100100110110000000000001000111000111110000000000000000000111100111110000000000000000000111000011110000000000000000000011000000110000000000000000000011000100110000000000000000000010011010110000000000000000000010011010110110000000000000000010011010110000000000000001000010011010110110000000000001000110011011110000000000000000000010000010110000000000000001000010000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam hphy_inst.m_hphy_ac_rom_init_file = "hps_ac_rom.hex";
defparam hphy_inst.m_hphy_inst_rom_content = 2560'b1000000000000000000010000000011010000000000010000001100000000000100000100000000000001000001010000000000010000011000000000000100000111000000000001000000100000000000010000100100000000000100001010000000000001000010110000000000010000110000000000000100001000000000000000000100000000000000010000110100000000000000010001000000000001010011010000000100000000110100000000000000010010000000010000000011010000000000000001001100000000000101001101000000000001000011010000000100000000110100000000000000010110110100000001100110011101000000000001010111010000000100011001110100000000000101110001000000011101100100010000000000010100000100000001010110010001000100000000110100000000000110011100000000000001100110110000000000011100111000000000000000011000000000000100000110011100000001000001100111000000010000011001110000000100000110011100000000000001101000000000000000001101000000000000000011010000000000000000110100000000000000001101000000001100000111010000000011000010000100000000110000100001000000001100001000010000000000010100110100000000000100001101000000010000000011010000000000011001110000000000000110011011000000000001110011100000000000000001100000000000011000011001110000000110000110011100000001100001100111000000011000011001110000000000000110100000000000000000110100000000000000001101000000000000000011010000000000000000110100000000111000011101000000001110001000010000000011100010000100000000111000100001000000000001010011010000000000010000110100000001000000001101000000000000001000101011000000000000110110110001000000001101000000000000001000101101000000000000111111010000000000001111110100000001000011111101000010000001111111010000100000100001110100001000001000011101000010000010000111010000000000100010110100000000000011111101000000000000111111010000000101001111110100010000000011010000000010000001110100010000100000100001000100001000001000010001000010000010000100010000100000011110110100001000001000011101000010000010000111010000100000100001110100000001010011010000000010000001111111010000100000100001110100001000001000011101000010000010000111010000100000100000000100001000001000010001000010000010000100010000100000100001000100000000001000100000000000011000110100000000000100001101000000000001110011010000000100000000110100000000000000000000000000000001000000000000000000010100000000000000000110000000000000010000000000000000000000000000000100000000000100000001000000000001010000010000000000011000000100000001000000000001000000000001001000110000000000010000110100000000000101001101000000010000000011010000000010000001111000010001000000001101000000000000000000000000000;
defparam hphy_inst.m_hphy_inst_rom_init_file = "hps_inst_rom.hex";

endmodule

module terminal_qsys_hps_sdram_p0_acv_hard_io_pads (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	dqsin1,
	pad_gen0raw_input1,
	pad_gen1raw_input1,
	pad_gen2raw_input1,
	pad_gen3raw_input1,
	pad_gen4raw_input1,
	pad_gen5raw_input1,
	pad_gen6raw_input1,
	pad_gen7raw_input1,
	dqsin2,
	pad_gen0raw_input2,
	pad_gen1raw_input2,
	pad_gen2raw_input2,
	pad_gen3raw_input2,
	pad_gen4raw_input2,
	pad_gen5raw_input2,
	pad_gen6raw_input2,
	pad_gen7raw_input2,
	dqsin3,
	pad_gen0raw_input3,
	pad_gen1raw_input3,
	pad_gen2raw_input3,
	pad_gen3raw_input3,
	pad_gen4raw_input3,
	pad_gen5raw_input3,
	pad_gen6raw_input3,
	pad_gen7raw_input3,
	afi_clk,
	pll_write_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	extra_output_pad_gen0delayed_data_out,
	extra_output_pad_gen0delayed_data_out1,
	extra_output_pad_gen0delayed_data_out2,
	extra_output_pad_gen0delayed_data_out3,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	pad_gen0delayed_data_out1,
	pad_gen0delayed_oe_11,
	delayed_oct1,
	pad_gen1delayed_data_out1,
	pad_gen1delayed_oe_11,
	pad_gen2delayed_data_out1,
	pad_gen2delayed_oe_11,
	pad_gen3delayed_data_out1,
	pad_gen3delayed_oe_11,
	pad_gen4delayed_data_out1,
	pad_gen4delayed_oe_11,
	pad_gen5delayed_data_out1,
	pad_gen5delayed_oe_11,
	pad_gen6delayed_data_out1,
	pad_gen6delayed_oe_11,
	pad_gen7delayed_data_out1,
	pad_gen7delayed_oe_11,
	pad_gen0delayed_data_out2,
	pad_gen0delayed_oe_12,
	delayed_oct2,
	pad_gen1delayed_data_out2,
	pad_gen1delayed_oe_12,
	pad_gen2delayed_data_out2,
	pad_gen2delayed_oe_12,
	pad_gen3delayed_data_out2,
	pad_gen3delayed_oe_12,
	pad_gen4delayed_data_out2,
	pad_gen4delayed_oe_12,
	pad_gen5delayed_data_out2,
	pad_gen5delayed_oe_12,
	pad_gen6delayed_data_out2,
	pad_gen6delayed_oe_12,
	pad_gen7delayed_data_out2,
	pad_gen7delayed_oe_12,
	pad_gen0delayed_data_out3,
	pad_gen0delayed_oe_13,
	delayed_oct3,
	pad_gen1delayed_data_out3,
	pad_gen1delayed_oe_13,
	pad_gen2delayed_data_out3,
	pad_gen2delayed_oe_13,
	pad_gen3delayed_data_out3,
	pad_gen3delayed_oe_13,
	pad_gen4delayed_data_out3,
	pad_gen4delayed_oe_13,
	pad_gen5delayed_data_out3,
	pad_gen5delayed_oe_13,
	pad_gen6delayed_data_out3,
	pad_gen6delayed_oe_13,
	pad_gen7delayed_data_out3,
	pad_gen7delayed_oe_13,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	os1,
	os_bar1,
	diff_oe1,
	diff_oe_bar1,
	diff_dtc1,
	diff_dtc_bar1,
	os2,
	os_bar2,
	diff_oe2,
	diff_oe_bar2,
	diff_dtc2,
	diff_dtc_bar2,
	os3,
	os_bar3,
	diff_oe3,
	diff_oe_bar3,
	diff_dtc3,
	diff_dtc_bar3,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	input_path_gen0read_fifo_out_01,
	input_path_gen0read_fifo_out_11,
	input_path_gen0read_fifo_out_21,
	input_path_gen0read_fifo_out_31,
	input_path_gen1read_fifo_out_01,
	input_path_gen1read_fifo_out_11,
	input_path_gen1read_fifo_out_21,
	input_path_gen1read_fifo_out_31,
	input_path_gen2read_fifo_out_01,
	input_path_gen2read_fifo_out_11,
	input_path_gen2read_fifo_out_21,
	input_path_gen2read_fifo_out_31,
	input_path_gen3read_fifo_out_01,
	input_path_gen3read_fifo_out_11,
	input_path_gen3read_fifo_out_21,
	input_path_gen3read_fifo_out_31,
	input_path_gen4read_fifo_out_01,
	input_path_gen4read_fifo_out_11,
	input_path_gen4read_fifo_out_21,
	input_path_gen4read_fifo_out_31,
	input_path_gen5read_fifo_out_01,
	input_path_gen5read_fifo_out_11,
	input_path_gen5read_fifo_out_21,
	input_path_gen5read_fifo_out_31,
	input_path_gen6read_fifo_out_01,
	input_path_gen6read_fifo_out_11,
	input_path_gen6read_fifo_out_21,
	input_path_gen6read_fifo_out_31,
	input_path_gen7read_fifo_out_01,
	input_path_gen7read_fifo_out_11,
	input_path_gen7read_fifo_out_21,
	input_path_gen7read_fifo_out_31,
	input_path_gen0read_fifo_out_02,
	input_path_gen0read_fifo_out_12,
	input_path_gen0read_fifo_out_22,
	input_path_gen0read_fifo_out_32,
	input_path_gen1read_fifo_out_02,
	input_path_gen1read_fifo_out_12,
	input_path_gen1read_fifo_out_22,
	input_path_gen1read_fifo_out_32,
	input_path_gen2read_fifo_out_02,
	input_path_gen2read_fifo_out_12,
	input_path_gen2read_fifo_out_22,
	input_path_gen2read_fifo_out_32,
	input_path_gen3read_fifo_out_02,
	input_path_gen3read_fifo_out_12,
	input_path_gen3read_fifo_out_22,
	input_path_gen3read_fifo_out_32,
	input_path_gen4read_fifo_out_02,
	input_path_gen4read_fifo_out_12,
	input_path_gen4read_fifo_out_22,
	input_path_gen4read_fifo_out_32,
	input_path_gen5read_fifo_out_02,
	input_path_gen5read_fifo_out_12,
	input_path_gen5read_fifo_out_22,
	input_path_gen5read_fifo_out_32,
	input_path_gen6read_fifo_out_02,
	input_path_gen6read_fifo_out_12,
	input_path_gen6read_fifo_out_22,
	input_path_gen6read_fifo_out_32,
	input_path_gen7read_fifo_out_02,
	input_path_gen7read_fifo_out_12,
	input_path_gen7read_fifo_out_22,
	input_path_gen7read_fifo_out_32,
	input_path_gen0read_fifo_out_03,
	input_path_gen0read_fifo_out_13,
	input_path_gen0read_fifo_out_23,
	input_path_gen0read_fifo_out_33,
	input_path_gen1read_fifo_out_03,
	input_path_gen1read_fifo_out_13,
	input_path_gen1read_fifo_out_23,
	input_path_gen1read_fifo_out_33,
	input_path_gen2read_fifo_out_03,
	input_path_gen2read_fifo_out_13,
	input_path_gen2read_fifo_out_23,
	input_path_gen2read_fifo_out_33,
	input_path_gen3read_fifo_out_03,
	input_path_gen3read_fifo_out_13,
	input_path_gen3read_fifo_out_23,
	input_path_gen3read_fifo_out_33,
	input_path_gen4read_fifo_out_03,
	input_path_gen4read_fifo_out_13,
	input_path_gen4read_fifo_out_23,
	input_path_gen4read_fifo_out_33,
	input_path_gen5read_fifo_out_03,
	input_path_gen5read_fifo_out_13,
	input_path_gen5read_fifo_out_23,
	input_path_gen5read_fifo_out_33,
	input_path_gen6read_fifo_out_03,
	input_path_gen6read_fifo_out_13,
	input_path_gen6read_fifo_out_23,
	input_path_gen6read_fifo_out_33,
	input_path_gen7read_fifo_out_03,
	input_path_gen7read_fifo_out_13,
	input_path_gen7read_fifo_out_23,
	input_path_gen7read_fifo_out_33,
	ddio_phy_dqslogic_rdatavalid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	dqsin1;
input 	pad_gen0raw_input1;
input 	pad_gen1raw_input1;
input 	pad_gen2raw_input1;
input 	pad_gen3raw_input1;
input 	pad_gen4raw_input1;
input 	pad_gen5raw_input1;
input 	pad_gen6raw_input1;
input 	pad_gen7raw_input1;
input 	dqsin2;
input 	pad_gen0raw_input2;
input 	pad_gen1raw_input2;
input 	pad_gen2raw_input2;
input 	pad_gen3raw_input2;
input 	pad_gen4raw_input2;
input 	pad_gen5raw_input2;
input 	pad_gen6raw_input2;
input 	pad_gen7raw_input2;
input 	dqsin3;
input 	pad_gen0raw_input3;
input 	pad_gen1raw_input3;
input 	pad_gen2raw_input3;
input 	pad_gen3raw_input3;
input 	pad_gen4raw_input3;
input 	pad_gen5raw_input3;
input 	pad_gen6raw_input3;
input 	pad_gen7raw_input3;
input 	afi_clk;
input 	pll_write_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	extra_output_pad_gen0delayed_data_out;
output 	extra_output_pad_gen0delayed_data_out1;
output 	extra_output_pad_gen0delayed_data_out2;
output 	extra_output_pad_gen0delayed_data_out3;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	pad_gen0delayed_data_out1;
output 	pad_gen0delayed_oe_11;
output 	delayed_oct1;
output 	pad_gen1delayed_data_out1;
output 	pad_gen1delayed_oe_11;
output 	pad_gen2delayed_data_out1;
output 	pad_gen2delayed_oe_11;
output 	pad_gen3delayed_data_out1;
output 	pad_gen3delayed_oe_11;
output 	pad_gen4delayed_data_out1;
output 	pad_gen4delayed_oe_11;
output 	pad_gen5delayed_data_out1;
output 	pad_gen5delayed_oe_11;
output 	pad_gen6delayed_data_out1;
output 	pad_gen6delayed_oe_11;
output 	pad_gen7delayed_data_out1;
output 	pad_gen7delayed_oe_11;
output 	pad_gen0delayed_data_out2;
output 	pad_gen0delayed_oe_12;
output 	delayed_oct2;
output 	pad_gen1delayed_data_out2;
output 	pad_gen1delayed_oe_12;
output 	pad_gen2delayed_data_out2;
output 	pad_gen2delayed_oe_12;
output 	pad_gen3delayed_data_out2;
output 	pad_gen3delayed_oe_12;
output 	pad_gen4delayed_data_out2;
output 	pad_gen4delayed_oe_12;
output 	pad_gen5delayed_data_out2;
output 	pad_gen5delayed_oe_12;
output 	pad_gen6delayed_data_out2;
output 	pad_gen6delayed_oe_12;
output 	pad_gen7delayed_data_out2;
output 	pad_gen7delayed_oe_12;
output 	pad_gen0delayed_data_out3;
output 	pad_gen0delayed_oe_13;
output 	delayed_oct3;
output 	pad_gen1delayed_data_out3;
output 	pad_gen1delayed_oe_13;
output 	pad_gen2delayed_data_out3;
output 	pad_gen2delayed_oe_13;
output 	pad_gen3delayed_data_out3;
output 	pad_gen3delayed_oe_13;
output 	pad_gen4delayed_data_out3;
output 	pad_gen4delayed_oe_13;
output 	pad_gen5delayed_data_out3;
output 	pad_gen5delayed_oe_13;
output 	pad_gen6delayed_data_out3;
output 	pad_gen6delayed_oe_13;
output 	pad_gen7delayed_data_out3;
output 	pad_gen7delayed_oe_13;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	os1;
output 	os_bar1;
output 	diff_oe1;
output 	diff_oe_bar1;
output 	diff_dtc1;
output 	diff_dtc_bar1;
output 	os2;
output 	os_bar2;
output 	diff_oe2;
output 	diff_oe_bar2;
output 	diff_dtc2;
output 	diff_dtc_bar2;
output 	os3;
output 	os_bar3;
output 	diff_oe3;
output 	diff_oe_bar3;
output 	diff_dtc3;
output 	diff_dtc_bar3;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	input_path_gen0read_fifo_out_01;
output 	input_path_gen0read_fifo_out_11;
output 	input_path_gen0read_fifo_out_21;
output 	input_path_gen0read_fifo_out_31;
output 	input_path_gen1read_fifo_out_01;
output 	input_path_gen1read_fifo_out_11;
output 	input_path_gen1read_fifo_out_21;
output 	input_path_gen1read_fifo_out_31;
output 	input_path_gen2read_fifo_out_01;
output 	input_path_gen2read_fifo_out_11;
output 	input_path_gen2read_fifo_out_21;
output 	input_path_gen2read_fifo_out_31;
output 	input_path_gen3read_fifo_out_01;
output 	input_path_gen3read_fifo_out_11;
output 	input_path_gen3read_fifo_out_21;
output 	input_path_gen3read_fifo_out_31;
output 	input_path_gen4read_fifo_out_01;
output 	input_path_gen4read_fifo_out_11;
output 	input_path_gen4read_fifo_out_21;
output 	input_path_gen4read_fifo_out_31;
output 	input_path_gen5read_fifo_out_01;
output 	input_path_gen5read_fifo_out_11;
output 	input_path_gen5read_fifo_out_21;
output 	input_path_gen5read_fifo_out_31;
output 	input_path_gen6read_fifo_out_01;
output 	input_path_gen6read_fifo_out_11;
output 	input_path_gen6read_fifo_out_21;
output 	input_path_gen6read_fifo_out_31;
output 	input_path_gen7read_fifo_out_01;
output 	input_path_gen7read_fifo_out_11;
output 	input_path_gen7read_fifo_out_21;
output 	input_path_gen7read_fifo_out_31;
output 	input_path_gen0read_fifo_out_02;
output 	input_path_gen0read_fifo_out_12;
output 	input_path_gen0read_fifo_out_22;
output 	input_path_gen0read_fifo_out_32;
output 	input_path_gen1read_fifo_out_02;
output 	input_path_gen1read_fifo_out_12;
output 	input_path_gen1read_fifo_out_22;
output 	input_path_gen1read_fifo_out_32;
output 	input_path_gen2read_fifo_out_02;
output 	input_path_gen2read_fifo_out_12;
output 	input_path_gen2read_fifo_out_22;
output 	input_path_gen2read_fifo_out_32;
output 	input_path_gen3read_fifo_out_02;
output 	input_path_gen3read_fifo_out_12;
output 	input_path_gen3read_fifo_out_22;
output 	input_path_gen3read_fifo_out_32;
output 	input_path_gen4read_fifo_out_02;
output 	input_path_gen4read_fifo_out_12;
output 	input_path_gen4read_fifo_out_22;
output 	input_path_gen4read_fifo_out_32;
output 	input_path_gen5read_fifo_out_02;
output 	input_path_gen5read_fifo_out_12;
output 	input_path_gen5read_fifo_out_22;
output 	input_path_gen5read_fifo_out_32;
output 	input_path_gen6read_fifo_out_02;
output 	input_path_gen6read_fifo_out_12;
output 	input_path_gen6read_fifo_out_22;
output 	input_path_gen6read_fifo_out_32;
output 	input_path_gen7read_fifo_out_02;
output 	input_path_gen7read_fifo_out_12;
output 	input_path_gen7read_fifo_out_22;
output 	input_path_gen7read_fifo_out_32;
output 	input_path_gen0read_fifo_out_03;
output 	input_path_gen0read_fifo_out_13;
output 	input_path_gen0read_fifo_out_23;
output 	input_path_gen0read_fifo_out_33;
output 	input_path_gen1read_fifo_out_03;
output 	input_path_gen1read_fifo_out_13;
output 	input_path_gen1read_fifo_out_23;
output 	input_path_gen1read_fifo_out_33;
output 	input_path_gen2read_fifo_out_03;
output 	input_path_gen2read_fifo_out_13;
output 	input_path_gen2read_fifo_out_23;
output 	input_path_gen2read_fifo_out_33;
output 	input_path_gen3read_fifo_out_03;
output 	input_path_gen3read_fifo_out_13;
output 	input_path_gen3read_fifo_out_23;
output 	input_path_gen3read_fifo_out_33;
output 	input_path_gen4read_fifo_out_03;
output 	input_path_gen4read_fifo_out_13;
output 	input_path_gen4read_fifo_out_23;
output 	input_path_gen4read_fifo_out_33;
output 	input_path_gen5read_fifo_out_03;
output 	input_path_gen5read_fifo_out_13;
output 	input_path_gen5read_fifo_out_23;
output 	input_path_gen5read_fifo_out_33;
output 	input_path_gen6read_fifo_out_03;
output 	input_path_gen6read_fifo_out_13;
output 	input_path_gen6read_fifo_out_23;
output 	input_path_gen6read_fifo_out_33;
output 	input_path_gen7read_fifo_out_03;
output 	input_path_gen7read_fifo_out_13;
output 	input_path_gen7read_fifo_out_23;
output 	input_path_gen7read_fifo_out_33;
output 	[4:0] ddio_phy_dqslogic_rdatavalid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_hps_sdram_p0_acv_hard_addr_cmd_pads uaddr_cmd_pads(
	.afi_clk(afi_clk),
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.dataout_9(dataout_9),
	.dataout_10(dataout_10),
	.dataout_11(dataout_11),
	.dataout_12(dataout_12),
	.dataout_13(dataout_13),
	.dataout_14(dataout_14),
	.dataout_01(dataout_01),
	.dataout_15(dataout_15),
	.dataout_21(dataout_21),
	.dataout_16(dataout_16),
	.dataout_02(dataout_02),
	.dataout_31(dataout_31),
	.dataout_41(dataout_41),
	.dataout_51(dataout_51),
	.dataout_03(dataout_03),
	.dataout_22(dataout_22),
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.phy_ddio_address_0(phy_ddio_address_0),
	.phy_ddio_address_1(phy_ddio_address_1),
	.phy_ddio_address_2(phy_ddio_address_2),
	.phy_ddio_address_3(phy_ddio_address_3),
	.phy_ddio_address_4(phy_ddio_address_4),
	.phy_ddio_address_5(phy_ddio_address_5),
	.phy_ddio_address_6(phy_ddio_address_6),
	.phy_ddio_address_7(phy_ddio_address_7),
	.phy_ddio_address_8(phy_ddio_address_8),
	.phy_ddio_address_9(phy_ddio_address_9),
	.phy_ddio_address_10(phy_ddio_address_10),
	.phy_ddio_address_11(phy_ddio_address_11),
	.phy_ddio_address_12(phy_ddio_address_12),
	.phy_ddio_address_13(phy_ddio_address_13),
	.phy_ddio_address_14(phy_ddio_address_14),
	.phy_ddio_address_15(phy_ddio_address_15),
	.phy_ddio_address_16(phy_ddio_address_16),
	.phy_ddio_address_17(phy_ddio_address_17),
	.phy_ddio_address_18(phy_ddio_address_18),
	.phy_ddio_address_19(phy_ddio_address_19),
	.phy_ddio_address_20(phy_ddio_address_20),
	.phy_ddio_address_21(phy_ddio_address_21),
	.phy_ddio_address_22(phy_ddio_address_22),
	.phy_ddio_address_23(phy_ddio_address_23),
	.phy_ddio_address_24(phy_ddio_address_24),
	.phy_ddio_address_25(phy_ddio_address_25),
	.phy_ddio_address_26(phy_ddio_address_26),
	.phy_ddio_address_27(phy_ddio_address_27),
	.phy_ddio_address_28(phy_ddio_address_28),
	.phy_ddio_address_29(phy_ddio_address_29),
	.phy_ddio_address_30(phy_ddio_address_30),
	.phy_ddio_address_31(phy_ddio_address_31),
	.phy_ddio_address_32(phy_ddio_address_32),
	.phy_ddio_address_33(phy_ddio_address_33),
	.phy_ddio_address_34(phy_ddio_address_34),
	.phy_ddio_address_35(phy_ddio_address_35),
	.phy_ddio_address_36(phy_ddio_address_36),
	.phy_ddio_address_37(phy_ddio_address_37),
	.phy_ddio_address_38(phy_ddio_address_38),
	.phy_ddio_address_39(phy_ddio_address_39),
	.phy_ddio_address_40(phy_ddio_address_40),
	.phy_ddio_address_41(phy_ddio_address_41),
	.phy_ddio_address_42(phy_ddio_address_42),
	.phy_ddio_address_43(phy_ddio_address_43),
	.phy_ddio_address_44(phy_ddio_address_44),
	.phy_ddio_address_45(phy_ddio_address_45),
	.phy_ddio_address_46(phy_ddio_address_46),
	.phy_ddio_address_47(phy_ddio_address_47),
	.phy_ddio_address_48(phy_ddio_address_48),
	.phy_ddio_address_49(phy_ddio_address_49),
	.phy_ddio_address_50(phy_ddio_address_50),
	.phy_ddio_address_51(phy_ddio_address_51),
	.phy_ddio_address_52(phy_ddio_address_52),
	.phy_ddio_address_53(phy_ddio_address_53),
	.phy_ddio_address_54(phy_ddio_address_54),
	.phy_ddio_address_55(phy_ddio_address_55),
	.phy_ddio_address_56(phy_ddio_address_56),
	.phy_ddio_address_57(phy_ddio_address_57),
	.phy_ddio_address_58(phy_ddio_address_58),
	.phy_ddio_address_59(phy_ddio_address_59),
	.phy_ddio_bank_0(phy_ddio_bank_0),
	.phy_ddio_bank_1(phy_ddio_bank_1),
	.phy_ddio_bank_2(phy_ddio_bank_2),
	.phy_ddio_bank_3(phy_ddio_bank_3),
	.phy_ddio_bank_4(phy_ddio_bank_4),
	.phy_ddio_bank_5(phy_ddio_bank_5),
	.phy_ddio_bank_6(phy_ddio_bank_6),
	.phy_ddio_bank_7(phy_ddio_bank_7),
	.phy_ddio_bank_8(phy_ddio_bank_8),
	.phy_ddio_bank_9(phy_ddio_bank_9),
	.phy_ddio_bank_10(phy_ddio_bank_10),
	.phy_ddio_bank_11(phy_ddio_bank_11),
	.phy_ddio_cas_n_0(phy_ddio_cas_n_0),
	.phy_ddio_cas_n_1(phy_ddio_cas_n_1),
	.phy_ddio_cas_n_2(phy_ddio_cas_n_2),
	.phy_ddio_cas_n_3(phy_ddio_cas_n_3),
	.phy_ddio_ck_0(phy_ddio_ck_0),
	.phy_ddio_ck_1(phy_ddio_ck_1),
	.phy_ddio_cke_0(phy_ddio_cke_0),
	.phy_ddio_cke_1(phy_ddio_cke_1),
	.phy_ddio_cke_2(phy_ddio_cke_2),
	.phy_ddio_cke_3(phy_ddio_cke_3),
	.phy_ddio_cs_n_0(phy_ddio_cs_n_0),
	.phy_ddio_cs_n_1(phy_ddio_cs_n_1),
	.phy_ddio_cs_n_2(phy_ddio_cs_n_2),
	.phy_ddio_cs_n_3(phy_ddio_cs_n_3),
	.phy_ddio_odt_0(phy_ddio_odt_0),
	.phy_ddio_odt_1(phy_ddio_odt_1),
	.phy_ddio_odt_2(phy_ddio_odt_2),
	.phy_ddio_odt_3(phy_ddio_odt_3),
	.phy_ddio_ras_n_0(phy_ddio_ras_n_0),
	.phy_ddio_ras_n_1(phy_ddio_ras_n_1),
	.phy_ddio_ras_n_2(phy_ddio_ras_n_2),
	.phy_ddio_ras_n_3(phy_ddio_ras_n_3),
	.phy_ddio_reset_n_0(phy_ddio_reset_n_0),
	.phy_ddio_reset_n_1(phy_ddio_reset_n_1),
	.phy_ddio_reset_n_2(phy_ddio_reset_n_2),
	.phy_ddio_reset_n_3(phy_ddio_reset_n_3),
	.phy_ddio_we_n_0(phy_ddio_we_n_0),
	.phy_ddio_we_n_1(phy_ddio_we_n_1),
	.phy_ddio_we_n_2(phy_ddio_we_n_2),
	.phy_ddio_we_n_3(phy_ddio_we_n_3),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6));

terminal_qsys_hps_sdram_p0_altdqdqs \dq_ddio[0].ubidir_dq_dqs (
	.dqsin(dqsin3),
	.pad_gen0raw_input(pad_gen0raw_input3),
	.pad_gen1raw_input(pad_gen1raw_input3),
	.pad_gen2raw_input(pad_gen2raw_input3),
	.pad_gen3raw_input(pad_gen3raw_input3),
	.pad_gen4raw_input(pad_gen4raw_input3),
	.pad_gen5raw_input(pad_gen5raw_input3),
	.pad_gen6raw_input(pad_gen6raw_input3),
	.pad_gen7raw_input(pad_gen7raw_input3),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out3),
	.phy_ddio_dmdout_0(phy_ddio_dmdout_0),
	.phy_ddio_dmdout_1(phy_ddio_dmdout_1),
	.phy_ddio_dmdout_2(phy_ddio_dmdout_2),
	.phy_ddio_dmdout_3(phy_ddio_dmdout_3),
	.phy_ddio_dqdout_0(phy_ddio_dqdout_0),
	.phy_ddio_dqdout_1(phy_ddio_dqdout_1),
	.phy_ddio_dqdout_2(phy_ddio_dqdout_2),
	.phy_ddio_dqdout_3(phy_ddio_dqdout_3),
	.phy_ddio_dqdout_4(phy_ddio_dqdout_4),
	.phy_ddio_dqdout_5(phy_ddio_dqdout_5),
	.phy_ddio_dqdout_6(phy_ddio_dqdout_6),
	.phy_ddio_dqdout_7(phy_ddio_dqdout_7),
	.phy_ddio_dqdout_8(phy_ddio_dqdout_8),
	.phy_ddio_dqdout_9(phy_ddio_dqdout_9),
	.phy_ddio_dqdout_10(phy_ddio_dqdout_10),
	.phy_ddio_dqdout_11(phy_ddio_dqdout_11),
	.phy_ddio_dqdout_12(phy_ddio_dqdout_12),
	.phy_ddio_dqdout_13(phy_ddio_dqdout_13),
	.phy_ddio_dqdout_14(phy_ddio_dqdout_14),
	.phy_ddio_dqdout_15(phy_ddio_dqdout_15),
	.phy_ddio_dqdout_16(phy_ddio_dqdout_16),
	.phy_ddio_dqdout_17(phy_ddio_dqdout_17),
	.phy_ddio_dqdout_18(phy_ddio_dqdout_18),
	.phy_ddio_dqdout_19(phy_ddio_dqdout_19),
	.phy_ddio_dqdout_20(phy_ddio_dqdout_20),
	.phy_ddio_dqdout_21(phy_ddio_dqdout_21),
	.phy_ddio_dqdout_22(phy_ddio_dqdout_22),
	.phy_ddio_dqdout_23(phy_ddio_dqdout_23),
	.phy_ddio_dqdout_24(phy_ddio_dqdout_24),
	.phy_ddio_dqdout_25(phy_ddio_dqdout_25),
	.phy_ddio_dqdout_26(phy_ddio_dqdout_26),
	.phy_ddio_dqdout_27(phy_ddio_dqdout_27),
	.phy_ddio_dqdout_28(phy_ddio_dqdout_28),
	.phy_ddio_dqdout_29(phy_ddio_dqdout_29),
	.phy_ddio_dqdout_30(phy_ddio_dqdout_30),
	.phy_ddio_dqdout_31(phy_ddio_dqdout_31),
	.phy_ddio_dqoe_0(phy_ddio_dqoe_0),
	.phy_ddio_dqoe_1(phy_ddio_dqoe_1),
	.phy_ddio_dqoe_2(phy_ddio_dqoe_2),
	.phy_ddio_dqoe_3(phy_ddio_dqoe_3),
	.phy_ddio_dqoe_4(phy_ddio_dqoe_4),
	.phy_ddio_dqoe_5(phy_ddio_dqoe_5),
	.phy_ddio_dqoe_6(phy_ddio_dqoe_6),
	.phy_ddio_dqoe_7(phy_ddio_dqoe_7),
	.phy_ddio_dqoe_8(phy_ddio_dqoe_8),
	.phy_ddio_dqoe_9(phy_ddio_dqoe_9),
	.phy_ddio_dqoe_10(phy_ddio_dqoe_10),
	.phy_ddio_dqoe_11(phy_ddio_dqoe_11),
	.phy_ddio_dqoe_12(phy_ddio_dqoe_12),
	.phy_ddio_dqoe_13(phy_ddio_dqoe_13),
	.phy_ddio_dqoe_14(phy_ddio_dqoe_14),
	.phy_ddio_dqoe_15(phy_ddio_dqoe_15),
	.phy_ddio_dqs_dout_0(phy_ddio_dqs_dout_0),
	.phy_ddio_dqs_dout_1(phy_ddio_dqs_dout_1),
	.phy_ddio_dqs_dout_2(phy_ddio_dqs_dout_2),
	.phy_ddio_dqs_dout_3(phy_ddio_dqs_dout_3),
	.phy_ddio_dqslogic_aclr_fifoctrl_0(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.phy_ddio_dqslogic_aclr_pstamble_0(phy_ddio_dqslogic_aclr_pstamble_0),
	.phy_ddio_dqslogic_dqsena_0(phy_ddio_dqslogic_dqsena_0),
	.phy_ddio_dqslogic_dqsena_1(phy_ddio_dqslogic_dqsena_1),
	.phy_ddio_dqslogic_fiforeset_0(phy_ddio_dqslogic_fiforeset_0),
	.phy_ddio_dqslogic_incrdataen_0(phy_ddio_dqslogic_incrdataen_0),
	.phy_ddio_dqslogic_incrdataen_1(phy_ddio_dqslogic_incrdataen_1),
	.phy_ddio_dqslogic_incwrptr_0(phy_ddio_dqslogic_incwrptr_0),
	.phy_ddio_dqslogic_incwrptr_1(phy_ddio_dqslogic_incwrptr_1),
	.phy_ddio_dqslogic_oct_0(phy_ddio_dqslogic_oct_0),
	.phy_ddio_dqslogic_oct_1(phy_ddio_dqslogic_oct_1),
	.phy_ddio_dqslogic_readlatency_0(phy_ddio_dqslogic_readlatency_0),
	.phy_ddio_dqslogic_readlatency_1(phy_ddio_dqslogic_readlatency_1),
	.phy_ddio_dqslogic_readlatency_2(phy_ddio_dqslogic_readlatency_2),
	.phy_ddio_dqslogic_readlatency_3(phy_ddio_dqslogic_readlatency_3),
	.phy_ddio_dqslogic_readlatency_4(phy_ddio_dqslogic_readlatency_4),
	.phy_ddio_dqs_oe_0(phy_ddio_dqs_oe_0),
	.phy_ddio_dqs_oe_1(phy_ddio_dqs_oe_1),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_0),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_1),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_2),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_3),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_0),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_1),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_2),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_3),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_0),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_1),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_2),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_3),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_0),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_1),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_2),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_3),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_0),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_1),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_2),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_3),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_0),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_1),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_2),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_3),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_0),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_1),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_2),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_3),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_0),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_1),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_2),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_3),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[0]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

terminal_qsys_hps_sdram_p0_altdqdqs_3 \dq_ddio[3].ubidir_dq_dqs (
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.phy_ddio_dmdout_12(phy_ddio_dmdout_12),
	.phy_ddio_dmdout_13(phy_ddio_dmdout_13),
	.phy_ddio_dmdout_14(phy_ddio_dmdout_14),
	.phy_ddio_dmdout_15(phy_ddio_dmdout_15),
	.phy_ddio_dqdout_108(phy_ddio_dqdout_108),
	.phy_ddio_dqdout_109(phy_ddio_dqdout_109),
	.phy_ddio_dqdout_110(phy_ddio_dqdout_110),
	.phy_ddio_dqdout_111(phy_ddio_dqdout_111),
	.phy_ddio_dqdout_112(phy_ddio_dqdout_112),
	.phy_ddio_dqdout_113(phy_ddio_dqdout_113),
	.phy_ddio_dqdout_114(phy_ddio_dqdout_114),
	.phy_ddio_dqdout_115(phy_ddio_dqdout_115),
	.phy_ddio_dqdout_116(phy_ddio_dqdout_116),
	.phy_ddio_dqdout_117(phy_ddio_dqdout_117),
	.phy_ddio_dqdout_118(phy_ddio_dqdout_118),
	.phy_ddio_dqdout_119(phy_ddio_dqdout_119),
	.phy_ddio_dqdout_120(phy_ddio_dqdout_120),
	.phy_ddio_dqdout_121(phy_ddio_dqdout_121),
	.phy_ddio_dqdout_122(phy_ddio_dqdout_122),
	.phy_ddio_dqdout_123(phy_ddio_dqdout_123),
	.phy_ddio_dqdout_124(phy_ddio_dqdout_124),
	.phy_ddio_dqdout_125(phy_ddio_dqdout_125),
	.phy_ddio_dqdout_126(phy_ddio_dqdout_126),
	.phy_ddio_dqdout_127(phy_ddio_dqdout_127),
	.phy_ddio_dqdout_128(phy_ddio_dqdout_128),
	.phy_ddio_dqdout_129(phy_ddio_dqdout_129),
	.phy_ddio_dqdout_130(phy_ddio_dqdout_130),
	.phy_ddio_dqdout_131(phy_ddio_dqdout_131),
	.phy_ddio_dqdout_132(phy_ddio_dqdout_132),
	.phy_ddio_dqdout_133(phy_ddio_dqdout_133),
	.phy_ddio_dqdout_134(phy_ddio_dqdout_134),
	.phy_ddio_dqdout_135(phy_ddio_dqdout_135),
	.phy_ddio_dqdout_136(phy_ddio_dqdout_136),
	.phy_ddio_dqdout_137(phy_ddio_dqdout_137),
	.phy_ddio_dqdout_138(phy_ddio_dqdout_138),
	.phy_ddio_dqdout_139(phy_ddio_dqdout_139),
	.phy_ddio_dqoe_54(phy_ddio_dqoe_54),
	.phy_ddio_dqoe_55(phy_ddio_dqoe_55),
	.phy_ddio_dqoe_56(phy_ddio_dqoe_56),
	.phy_ddio_dqoe_57(phy_ddio_dqoe_57),
	.phy_ddio_dqoe_58(phy_ddio_dqoe_58),
	.phy_ddio_dqoe_59(phy_ddio_dqoe_59),
	.phy_ddio_dqoe_60(phy_ddio_dqoe_60),
	.phy_ddio_dqoe_61(phy_ddio_dqoe_61),
	.phy_ddio_dqoe_62(phy_ddio_dqoe_62),
	.phy_ddio_dqoe_63(phy_ddio_dqoe_63),
	.phy_ddio_dqoe_64(phy_ddio_dqoe_64),
	.phy_ddio_dqoe_65(phy_ddio_dqoe_65),
	.phy_ddio_dqoe_66(phy_ddio_dqoe_66),
	.phy_ddio_dqoe_67(phy_ddio_dqoe_67),
	.phy_ddio_dqoe_68(phy_ddio_dqoe_68),
	.phy_ddio_dqoe_69(phy_ddio_dqoe_69),
	.phy_ddio_dqs_dout_12(phy_ddio_dqs_dout_12),
	.phy_ddio_dqs_dout_13(phy_ddio_dqs_dout_13),
	.phy_ddio_dqs_dout_14(phy_ddio_dqs_dout_14),
	.phy_ddio_dqs_dout_15(phy_ddio_dqs_dout_15),
	.phy_ddio_dqslogic_aclr_fifoctrl_3(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.phy_ddio_dqslogic_aclr_pstamble_3(phy_ddio_dqslogic_aclr_pstamble_3),
	.phy_ddio_dqslogic_dqsena_6(phy_ddio_dqslogic_dqsena_6),
	.phy_ddio_dqslogic_dqsena_7(phy_ddio_dqslogic_dqsena_7),
	.phy_ddio_dqslogic_fiforeset_3(phy_ddio_dqslogic_fiforeset_3),
	.phy_ddio_dqslogic_incrdataen_6(phy_ddio_dqslogic_incrdataen_6),
	.phy_ddio_dqslogic_incrdataen_7(phy_ddio_dqslogic_incrdataen_7),
	.phy_ddio_dqslogic_incwrptr_6(phy_ddio_dqslogic_incwrptr_6),
	.phy_ddio_dqslogic_incwrptr_7(phy_ddio_dqslogic_incwrptr_7),
	.phy_ddio_dqslogic_oct_6(phy_ddio_dqslogic_oct_6),
	.phy_ddio_dqslogic_oct_7(phy_ddio_dqslogic_oct_7),
	.phy_ddio_dqslogic_readlatency_15(phy_ddio_dqslogic_readlatency_15),
	.phy_ddio_dqslogic_readlatency_16(phy_ddio_dqslogic_readlatency_16),
	.phy_ddio_dqslogic_readlatency_17(phy_ddio_dqslogic_readlatency_17),
	.phy_ddio_dqslogic_readlatency_18(phy_ddio_dqslogic_readlatency_18),
	.phy_ddio_dqslogic_readlatency_19(phy_ddio_dqslogic_readlatency_19),
	.phy_ddio_dqs_oe_6(phy_ddio_dqs_oe_6),
	.phy_ddio_dqs_oe_7(phy_ddio_dqs_oe_7),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out3),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_13),
	.delayed_oct(delayed_oct3),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out3),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_13),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out3),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_13),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out3),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_13),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out3),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_13),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out3),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_13),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out3),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_13),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out3),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_13),
	.os(os3),
	.os_bar(os_bar3),
	.diff_oe(diff_oe3),
	.diff_oe_bar(diff_oe_bar3),
	.diff_dtc(diff_dtc3),
	.diff_dtc_bar(diff_dtc_bar3),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_03),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_13),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_23),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_33),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_03),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_13),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_23),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_33),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_03),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_13),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_23),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_33),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_03),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_13),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_23),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_33),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_03),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_13),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_23),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_33),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_03),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_13),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_23),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_33),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_03),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_13),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_23),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_33),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_03),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_13),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_23),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_33),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[3]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

terminal_qsys_hps_sdram_p0_altdqdqs_2 \dq_ddio[2].ubidir_dq_dqs (
	.dqsin(dqsin1),
	.pad_gen0raw_input(pad_gen0raw_input1),
	.pad_gen1raw_input(pad_gen1raw_input1),
	.pad_gen2raw_input(pad_gen2raw_input1),
	.pad_gen3raw_input(pad_gen3raw_input1),
	.pad_gen4raw_input(pad_gen4raw_input1),
	.pad_gen5raw_input(pad_gen5raw_input1),
	.pad_gen6raw_input(pad_gen6raw_input1),
	.pad_gen7raw_input(pad_gen7raw_input1),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out1),
	.phy_ddio_dmdout_8(phy_ddio_dmdout_8),
	.phy_ddio_dmdout_9(phy_ddio_dmdout_9),
	.phy_ddio_dmdout_10(phy_ddio_dmdout_10),
	.phy_ddio_dmdout_11(phy_ddio_dmdout_11),
	.phy_ddio_dqdout_72(phy_ddio_dqdout_72),
	.phy_ddio_dqdout_73(phy_ddio_dqdout_73),
	.phy_ddio_dqdout_74(phy_ddio_dqdout_74),
	.phy_ddio_dqdout_75(phy_ddio_dqdout_75),
	.phy_ddio_dqdout_76(phy_ddio_dqdout_76),
	.phy_ddio_dqdout_77(phy_ddio_dqdout_77),
	.phy_ddio_dqdout_78(phy_ddio_dqdout_78),
	.phy_ddio_dqdout_79(phy_ddio_dqdout_79),
	.phy_ddio_dqdout_80(phy_ddio_dqdout_80),
	.phy_ddio_dqdout_81(phy_ddio_dqdout_81),
	.phy_ddio_dqdout_82(phy_ddio_dqdout_82),
	.phy_ddio_dqdout_83(phy_ddio_dqdout_83),
	.phy_ddio_dqdout_84(phy_ddio_dqdout_84),
	.phy_ddio_dqdout_85(phy_ddio_dqdout_85),
	.phy_ddio_dqdout_86(phy_ddio_dqdout_86),
	.phy_ddio_dqdout_87(phy_ddio_dqdout_87),
	.phy_ddio_dqdout_88(phy_ddio_dqdout_88),
	.phy_ddio_dqdout_89(phy_ddio_dqdout_89),
	.phy_ddio_dqdout_90(phy_ddio_dqdout_90),
	.phy_ddio_dqdout_91(phy_ddio_dqdout_91),
	.phy_ddio_dqdout_92(phy_ddio_dqdout_92),
	.phy_ddio_dqdout_93(phy_ddio_dqdout_93),
	.phy_ddio_dqdout_94(phy_ddio_dqdout_94),
	.phy_ddio_dqdout_95(phy_ddio_dqdout_95),
	.phy_ddio_dqdout_96(phy_ddio_dqdout_96),
	.phy_ddio_dqdout_97(phy_ddio_dqdout_97),
	.phy_ddio_dqdout_98(phy_ddio_dqdout_98),
	.phy_ddio_dqdout_99(phy_ddio_dqdout_99),
	.phy_ddio_dqdout_100(phy_ddio_dqdout_100),
	.phy_ddio_dqdout_101(phy_ddio_dqdout_101),
	.phy_ddio_dqdout_102(phy_ddio_dqdout_102),
	.phy_ddio_dqdout_103(phy_ddio_dqdout_103),
	.phy_ddio_dqoe_36(phy_ddio_dqoe_36),
	.phy_ddio_dqoe_37(phy_ddio_dqoe_37),
	.phy_ddio_dqoe_38(phy_ddio_dqoe_38),
	.phy_ddio_dqoe_39(phy_ddio_dqoe_39),
	.phy_ddio_dqoe_40(phy_ddio_dqoe_40),
	.phy_ddio_dqoe_41(phy_ddio_dqoe_41),
	.phy_ddio_dqoe_42(phy_ddio_dqoe_42),
	.phy_ddio_dqoe_43(phy_ddio_dqoe_43),
	.phy_ddio_dqoe_44(phy_ddio_dqoe_44),
	.phy_ddio_dqoe_45(phy_ddio_dqoe_45),
	.phy_ddio_dqoe_46(phy_ddio_dqoe_46),
	.phy_ddio_dqoe_47(phy_ddio_dqoe_47),
	.phy_ddio_dqoe_48(phy_ddio_dqoe_48),
	.phy_ddio_dqoe_49(phy_ddio_dqoe_49),
	.phy_ddio_dqoe_50(phy_ddio_dqoe_50),
	.phy_ddio_dqoe_51(phy_ddio_dqoe_51),
	.phy_ddio_dqs_dout_8(phy_ddio_dqs_dout_8),
	.phy_ddio_dqs_dout_9(phy_ddio_dqs_dout_9),
	.phy_ddio_dqs_dout_10(phy_ddio_dqs_dout_10),
	.phy_ddio_dqs_dout_11(phy_ddio_dqs_dout_11),
	.phy_ddio_dqslogic_aclr_fifoctrl_2(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.phy_ddio_dqslogic_aclr_pstamble_2(phy_ddio_dqslogic_aclr_pstamble_2),
	.phy_ddio_dqslogic_dqsena_4(phy_ddio_dqslogic_dqsena_4),
	.phy_ddio_dqslogic_dqsena_5(phy_ddio_dqslogic_dqsena_5),
	.phy_ddio_dqslogic_fiforeset_2(phy_ddio_dqslogic_fiforeset_2),
	.phy_ddio_dqslogic_incrdataen_4(phy_ddio_dqslogic_incrdataen_4),
	.phy_ddio_dqslogic_incrdataen_5(phy_ddio_dqslogic_incrdataen_5),
	.phy_ddio_dqslogic_incwrptr_4(phy_ddio_dqslogic_incwrptr_4),
	.phy_ddio_dqslogic_incwrptr_5(phy_ddio_dqslogic_incwrptr_5),
	.phy_ddio_dqslogic_oct_4(phy_ddio_dqslogic_oct_4),
	.phy_ddio_dqslogic_oct_5(phy_ddio_dqslogic_oct_5),
	.phy_ddio_dqslogic_readlatency_10(phy_ddio_dqslogic_readlatency_10),
	.phy_ddio_dqslogic_readlatency_11(phy_ddio_dqslogic_readlatency_11),
	.phy_ddio_dqslogic_readlatency_12(phy_ddio_dqslogic_readlatency_12),
	.phy_ddio_dqslogic_readlatency_13(phy_ddio_dqslogic_readlatency_13),
	.phy_ddio_dqslogic_readlatency_14(phy_ddio_dqslogic_readlatency_14),
	.phy_ddio_dqs_oe_4(phy_ddio_dqs_oe_4),
	.phy_ddio_dqs_oe_5(phy_ddio_dqs_oe_5),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out2),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_12),
	.delayed_oct(delayed_oct2),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out2),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_12),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out2),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_12),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out2),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_12),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out2),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_12),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out2),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_12),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out2),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_12),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out2),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_12),
	.os(os2),
	.os_bar(os_bar2),
	.diff_oe(diff_oe2),
	.diff_oe_bar(diff_oe_bar2),
	.diff_dtc(diff_dtc2),
	.diff_dtc_bar(diff_dtc_bar2),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_02),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_12),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_22),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_32),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_02),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_12),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_22),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_32),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_02),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_12),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_22),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_32),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_02),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_12),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_22),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_32),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_02),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_12),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_22),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_32),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_02),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_12),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_22),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_32),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_02),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_12),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_22),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_32),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_02),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_12),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_22),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_32),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[2]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

terminal_qsys_hps_sdram_p0_altdqdqs_1 \dq_ddio[1].ubidir_dq_dqs (
	.dqsin(dqsin2),
	.pad_gen0raw_input(pad_gen0raw_input2),
	.pad_gen1raw_input(pad_gen1raw_input2),
	.pad_gen2raw_input(pad_gen2raw_input2),
	.pad_gen3raw_input(pad_gen3raw_input2),
	.pad_gen4raw_input(pad_gen4raw_input2),
	.pad_gen5raw_input(pad_gen5raw_input2),
	.pad_gen6raw_input(pad_gen6raw_input2),
	.pad_gen7raw_input(pad_gen7raw_input2),
	.afi_clk(afi_clk),
	.pll_write_clk(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out2),
	.phy_ddio_dmdout_4(phy_ddio_dmdout_4),
	.phy_ddio_dmdout_5(phy_ddio_dmdout_5),
	.phy_ddio_dmdout_6(phy_ddio_dmdout_6),
	.phy_ddio_dmdout_7(phy_ddio_dmdout_7),
	.phy_ddio_dqdout_36(phy_ddio_dqdout_36),
	.phy_ddio_dqdout_37(phy_ddio_dqdout_37),
	.phy_ddio_dqdout_38(phy_ddio_dqdout_38),
	.phy_ddio_dqdout_39(phy_ddio_dqdout_39),
	.phy_ddio_dqdout_40(phy_ddio_dqdout_40),
	.phy_ddio_dqdout_41(phy_ddio_dqdout_41),
	.phy_ddio_dqdout_42(phy_ddio_dqdout_42),
	.phy_ddio_dqdout_43(phy_ddio_dqdout_43),
	.phy_ddio_dqdout_44(phy_ddio_dqdout_44),
	.phy_ddio_dqdout_45(phy_ddio_dqdout_45),
	.phy_ddio_dqdout_46(phy_ddio_dqdout_46),
	.phy_ddio_dqdout_47(phy_ddio_dqdout_47),
	.phy_ddio_dqdout_48(phy_ddio_dqdout_48),
	.phy_ddio_dqdout_49(phy_ddio_dqdout_49),
	.phy_ddio_dqdout_50(phy_ddio_dqdout_50),
	.phy_ddio_dqdout_51(phy_ddio_dqdout_51),
	.phy_ddio_dqdout_52(phy_ddio_dqdout_52),
	.phy_ddio_dqdout_53(phy_ddio_dqdout_53),
	.phy_ddio_dqdout_54(phy_ddio_dqdout_54),
	.phy_ddio_dqdout_55(phy_ddio_dqdout_55),
	.phy_ddio_dqdout_56(phy_ddio_dqdout_56),
	.phy_ddio_dqdout_57(phy_ddio_dqdout_57),
	.phy_ddio_dqdout_58(phy_ddio_dqdout_58),
	.phy_ddio_dqdout_59(phy_ddio_dqdout_59),
	.phy_ddio_dqdout_60(phy_ddio_dqdout_60),
	.phy_ddio_dqdout_61(phy_ddio_dqdout_61),
	.phy_ddio_dqdout_62(phy_ddio_dqdout_62),
	.phy_ddio_dqdout_63(phy_ddio_dqdout_63),
	.phy_ddio_dqdout_64(phy_ddio_dqdout_64),
	.phy_ddio_dqdout_65(phy_ddio_dqdout_65),
	.phy_ddio_dqdout_66(phy_ddio_dqdout_66),
	.phy_ddio_dqdout_67(phy_ddio_dqdout_67),
	.phy_ddio_dqoe_18(phy_ddio_dqoe_18),
	.phy_ddio_dqoe_19(phy_ddio_dqoe_19),
	.phy_ddio_dqoe_20(phy_ddio_dqoe_20),
	.phy_ddio_dqoe_21(phy_ddio_dqoe_21),
	.phy_ddio_dqoe_22(phy_ddio_dqoe_22),
	.phy_ddio_dqoe_23(phy_ddio_dqoe_23),
	.phy_ddio_dqoe_24(phy_ddio_dqoe_24),
	.phy_ddio_dqoe_25(phy_ddio_dqoe_25),
	.phy_ddio_dqoe_26(phy_ddio_dqoe_26),
	.phy_ddio_dqoe_27(phy_ddio_dqoe_27),
	.phy_ddio_dqoe_28(phy_ddio_dqoe_28),
	.phy_ddio_dqoe_29(phy_ddio_dqoe_29),
	.phy_ddio_dqoe_30(phy_ddio_dqoe_30),
	.phy_ddio_dqoe_31(phy_ddio_dqoe_31),
	.phy_ddio_dqoe_32(phy_ddio_dqoe_32),
	.phy_ddio_dqoe_33(phy_ddio_dqoe_33),
	.phy_ddio_dqs_dout_4(phy_ddio_dqs_dout_4),
	.phy_ddio_dqs_dout_5(phy_ddio_dqs_dout_5),
	.phy_ddio_dqs_dout_6(phy_ddio_dqs_dout_6),
	.phy_ddio_dqs_dout_7(phy_ddio_dqs_dout_7),
	.phy_ddio_dqslogic_aclr_fifoctrl_1(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.phy_ddio_dqslogic_aclr_pstamble_1(phy_ddio_dqslogic_aclr_pstamble_1),
	.phy_ddio_dqslogic_dqsena_2(phy_ddio_dqslogic_dqsena_2),
	.phy_ddio_dqslogic_dqsena_3(phy_ddio_dqslogic_dqsena_3),
	.phy_ddio_dqslogic_fiforeset_1(phy_ddio_dqslogic_fiforeset_1),
	.phy_ddio_dqslogic_incrdataen_2(phy_ddio_dqslogic_incrdataen_2),
	.phy_ddio_dqslogic_incrdataen_3(phy_ddio_dqslogic_incrdataen_3),
	.phy_ddio_dqslogic_incwrptr_2(phy_ddio_dqslogic_incwrptr_2),
	.phy_ddio_dqslogic_incwrptr_3(phy_ddio_dqslogic_incwrptr_3),
	.phy_ddio_dqslogic_oct_2(phy_ddio_dqslogic_oct_2),
	.phy_ddio_dqslogic_oct_3(phy_ddio_dqslogic_oct_3),
	.phy_ddio_dqslogic_readlatency_5(phy_ddio_dqslogic_readlatency_5),
	.phy_ddio_dqslogic_readlatency_6(phy_ddio_dqslogic_readlatency_6),
	.phy_ddio_dqslogic_readlatency_7(phy_ddio_dqslogic_readlatency_7),
	.phy_ddio_dqslogic_readlatency_8(phy_ddio_dqslogic_readlatency_8),
	.phy_ddio_dqslogic_readlatency_9(phy_ddio_dqslogic_readlatency_9),
	.phy_ddio_dqs_oe_2(phy_ddio_dqs_oe_2),
	.phy_ddio_dqs_oe_3(phy_ddio_dqs_oe_3),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out1),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_11),
	.delayed_oct(delayed_oct1),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out1),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_11),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out1),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_11),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out1),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_11),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out1),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_11),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out1),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_11),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out1),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_11),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out1),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_11),
	.os(os1),
	.os_bar(os_bar1),
	.diff_oe(diff_oe1),
	.diff_oe_bar(diff_oe_bar1),
	.diff_dtc(diff_dtc1),
	.diff_dtc_bar(diff_dtc_bar1),
	.input_path_gen0read_fifo_out_0(input_path_gen0read_fifo_out_01),
	.input_path_gen0read_fifo_out_1(input_path_gen0read_fifo_out_11),
	.input_path_gen0read_fifo_out_2(input_path_gen0read_fifo_out_21),
	.input_path_gen0read_fifo_out_3(input_path_gen0read_fifo_out_31),
	.input_path_gen1read_fifo_out_0(input_path_gen1read_fifo_out_01),
	.input_path_gen1read_fifo_out_1(input_path_gen1read_fifo_out_11),
	.input_path_gen1read_fifo_out_2(input_path_gen1read_fifo_out_21),
	.input_path_gen1read_fifo_out_3(input_path_gen1read_fifo_out_31),
	.input_path_gen2read_fifo_out_0(input_path_gen2read_fifo_out_01),
	.input_path_gen2read_fifo_out_1(input_path_gen2read_fifo_out_11),
	.input_path_gen2read_fifo_out_2(input_path_gen2read_fifo_out_21),
	.input_path_gen2read_fifo_out_3(input_path_gen2read_fifo_out_31),
	.input_path_gen3read_fifo_out_0(input_path_gen3read_fifo_out_01),
	.input_path_gen3read_fifo_out_1(input_path_gen3read_fifo_out_11),
	.input_path_gen3read_fifo_out_2(input_path_gen3read_fifo_out_21),
	.input_path_gen3read_fifo_out_3(input_path_gen3read_fifo_out_31),
	.input_path_gen4read_fifo_out_0(input_path_gen4read_fifo_out_01),
	.input_path_gen4read_fifo_out_1(input_path_gen4read_fifo_out_11),
	.input_path_gen4read_fifo_out_2(input_path_gen4read_fifo_out_21),
	.input_path_gen4read_fifo_out_3(input_path_gen4read_fifo_out_31),
	.input_path_gen5read_fifo_out_0(input_path_gen5read_fifo_out_01),
	.input_path_gen5read_fifo_out_1(input_path_gen5read_fifo_out_11),
	.input_path_gen5read_fifo_out_2(input_path_gen5read_fifo_out_21),
	.input_path_gen5read_fifo_out_3(input_path_gen5read_fifo_out_31),
	.input_path_gen6read_fifo_out_0(input_path_gen6read_fifo_out_01),
	.input_path_gen6read_fifo_out_1(input_path_gen6read_fifo_out_11),
	.input_path_gen6read_fifo_out_2(input_path_gen6read_fifo_out_21),
	.input_path_gen6read_fifo_out_3(input_path_gen6read_fifo_out_31),
	.input_path_gen7read_fifo_out_0(input_path_gen7read_fifo_out_01),
	.input_path_gen7read_fifo_out_1(input_path_gen7read_fifo_out_11),
	.input_path_gen7read_fifo_out_2(input_path_gen7read_fifo_out_21),
	.input_path_gen7read_fifo_out_3(input_path_gen7read_fifo_out_31),
	.lfifo_rdata_valid(ddio_phy_dqslogic_rdatavalid[1]),
	.dll_delayctrl_0(dll_delayctrl_0),
	.dll_delayctrl_1(dll_delayctrl_1),
	.dll_delayctrl_2(dll_delayctrl_2),
	.dll_delayctrl_3(dll_delayctrl_3),
	.dll_delayctrl_4(dll_delayctrl_4),
	.dll_delayctrl_5(dll_delayctrl_5),
	.dll_delayctrl_6(dll_delayctrl_6),
	.GND_port(GND_port));

endmodule

module terminal_qsys_hps_sdram_p0_acv_hard_addr_cmd_pads (
	afi_clk,
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	dataout_9,
	dataout_10,
	dataout_11,
	dataout_12,
	dataout_13,
	dataout_14,
	dataout_01,
	dataout_15,
	dataout_21,
	dataout_16,
	dataout_02,
	dataout_31,
	dataout_41,
	dataout_51,
	dataout_03,
	dataout_22,
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	phy_ddio_address_0,
	phy_ddio_address_1,
	phy_ddio_address_2,
	phy_ddio_address_3,
	phy_ddio_address_4,
	phy_ddio_address_5,
	phy_ddio_address_6,
	phy_ddio_address_7,
	phy_ddio_address_8,
	phy_ddio_address_9,
	phy_ddio_address_10,
	phy_ddio_address_11,
	phy_ddio_address_12,
	phy_ddio_address_13,
	phy_ddio_address_14,
	phy_ddio_address_15,
	phy_ddio_address_16,
	phy_ddio_address_17,
	phy_ddio_address_18,
	phy_ddio_address_19,
	phy_ddio_address_20,
	phy_ddio_address_21,
	phy_ddio_address_22,
	phy_ddio_address_23,
	phy_ddio_address_24,
	phy_ddio_address_25,
	phy_ddio_address_26,
	phy_ddio_address_27,
	phy_ddio_address_28,
	phy_ddio_address_29,
	phy_ddio_address_30,
	phy_ddio_address_31,
	phy_ddio_address_32,
	phy_ddio_address_33,
	phy_ddio_address_34,
	phy_ddio_address_35,
	phy_ddio_address_36,
	phy_ddio_address_37,
	phy_ddio_address_38,
	phy_ddio_address_39,
	phy_ddio_address_40,
	phy_ddio_address_41,
	phy_ddio_address_42,
	phy_ddio_address_43,
	phy_ddio_address_44,
	phy_ddio_address_45,
	phy_ddio_address_46,
	phy_ddio_address_47,
	phy_ddio_address_48,
	phy_ddio_address_49,
	phy_ddio_address_50,
	phy_ddio_address_51,
	phy_ddio_address_52,
	phy_ddio_address_53,
	phy_ddio_address_54,
	phy_ddio_address_55,
	phy_ddio_address_56,
	phy_ddio_address_57,
	phy_ddio_address_58,
	phy_ddio_address_59,
	phy_ddio_bank_0,
	phy_ddio_bank_1,
	phy_ddio_bank_2,
	phy_ddio_bank_3,
	phy_ddio_bank_4,
	phy_ddio_bank_5,
	phy_ddio_bank_6,
	phy_ddio_bank_7,
	phy_ddio_bank_8,
	phy_ddio_bank_9,
	phy_ddio_bank_10,
	phy_ddio_bank_11,
	phy_ddio_cas_n_0,
	phy_ddio_cas_n_1,
	phy_ddio_cas_n_2,
	phy_ddio_cas_n_3,
	phy_ddio_ck_0,
	phy_ddio_ck_1,
	phy_ddio_cke_0,
	phy_ddio_cke_1,
	phy_ddio_cke_2,
	phy_ddio_cke_3,
	phy_ddio_cs_n_0,
	phy_ddio_cs_n_1,
	phy_ddio_cs_n_2,
	phy_ddio_cs_n_3,
	phy_ddio_odt_0,
	phy_ddio_odt_1,
	phy_ddio_odt_2,
	phy_ddio_odt_3,
	phy_ddio_ras_n_0,
	phy_ddio_ras_n_1,
	phy_ddio_ras_n_2,
	phy_ddio_ras_n_3,
	phy_ddio_reset_n_0,
	phy_ddio_reset_n_1,
	phy_ddio_reset_n_2,
	phy_ddio_reset_n_3,
	phy_ddio_we_n_0,
	phy_ddio_we_n_1,
	phy_ddio_we_n_2,
	phy_ddio_we_n_3,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6)/* synthesis synthesis_greybox=0 */;
input 	afi_clk;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
output 	dataout_9;
output 	dataout_10;
output 	dataout_11;
output 	dataout_12;
output 	dataout_13;
output 	dataout_14;
output 	dataout_01;
output 	dataout_15;
output 	dataout_21;
output 	dataout_16;
output 	dataout_02;
output 	dataout_31;
output 	dataout_41;
output 	dataout_51;
output 	dataout_03;
output 	dataout_22;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	phy_ddio_address_0;
input 	phy_ddio_address_1;
input 	phy_ddio_address_2;
input 	phy_ddio_address_3;
input 	phy_ddio_address_4;
input 	phy_ddio_address_5;
input 	phy_ddio_address_6;
input 	phy_ddio_address_7;
input 	phy_ddio_address_8;
input 	phy_ddio_address_9;
input 	phy_ddio_address_10;
input 	phy_ddio_address_11;
input 	phy_ddio_address_12;
input 	phy_ddio_address_13;
input 	phy_ddio_address_14;
input 	phy_ddio_address_15;
input 	phy_ddio_address_16;
input 	phy_ddio_address_17;
input 	phy_ddio_address_18;
input 	phy_ddio_address_19;
input 	phy_ddio_address_20;
input 	phy_ddio_address_21;
input 	phy_ddio_address_22;
input 	phy_ddio_address_23;
input 	phy_ddio_address_24;
input 	phy_ddio_address_25;
input 	phy_ddio_address_26;
input 	phy_ddio_address_27;
input 	phy_ddio_address_28;
input 	phy_ddio_address_29;
input 	phy_ddio_address_30;
input 	phy_ddio_address_31;
input 	phy_ddio_address_32;
input 	phy_ddio_address_33;
input 	phy_ddio_address_34;
input 	phy_ddio_address_35;
input 	phy_ddio_address_36;
input 	phy_ddio_address_37;
input 	phy_ddio_address_38;
input 	phy_ddio_address_39;
input 	phy_ddio_address_40;
input 	phy_ddio_address_41;
input 	phy_ddio_address_42;
input 	phy_ddio_address_43;
input 	phy_ddio_address_44;
input 	phy_ddio_address_45;
input 	phy_ddio_address_46;
input 	phy_ddio_address_47;
input 	phy_ddio_address_48;
input 	phy_ddio_address_49;
input 	phy_ddio_address_50;
input 	phy_ddio_address_51;
input 	phy_ddio_address_52;
input 	phy_ddio_address_53;
input 	phy_ddio_address_54;
input 	phy_ddio_address_55;
input 	phy_ddio_address_56;
input 	phy_ddio_address_57;
input 	phy_ddio_address_58;
input 	phy_ddio_address_59;
input 	phy_ddio_bank_0;
input 	phy_ddio_bank_1;
input 	phy_ddio_bank_2;
input 	phy_ddio_bank_3;
input 	phy_ddio_bank_4;
input 	phy_ddio_bank_5;
input 	phy_ddio_bank_6;
input 	phy_ddio_bank_7;
input 	phy_ddio_bank_8;
input 	phy_ddio_bank_9;
input 	phy_ddio_bank_10;
input 	phy_ddio_bank_11;
input 	phy_ddio_cas_n_0;
input 	phy_ddio_cas_n_1;
input 	phy_ddio_cas_n_2;
input 	phy_ddio_cas_n_3;
input 	phy_ddio_ck_0;
input 	phy_ddio_ck_1;
input 	phy_ddio_cke_0;
input 	phy_ddio_cke_1;
input 	phy_ddio_cke_2;
input 	phy_ddio_cke_3;
input 	phy_ddio_cs_n_0;
input 	phy_ddio_cs_n_1;
input 	phy_ddio_cs_n_2;
input 	phy_ddio_cs_n_3;
input 	phy_ddio_odt_0;
input 	phy_ddio_odt_1;
input 	phy_ddio_odt_2;
input 	phy_ddio_odt_3;
input 	phy_ddio_ras_n_0;
input 	phy_ddio_ras_n_1;
input 	phy_ddio_ras_n_2;
input 	phy_ddio_ras_n_3;
input 	phy_ddio_reset_n_0;
input 	phy_ddio_reset_n_1;
input 	phy_ddio_reset_n_2;
input 	phy_ddio_reset_n_3;
input 	phy_ddio_we_n_0;
input 	phy_ddio_we_n_1;
input 	phy_ddio_we_n_2;
input 	phy_ddio_we_n_3;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_gen[0].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[1].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[2].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[3].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[4].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[5].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[6].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[7].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[8].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[9].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[10].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[11].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[12].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[13].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[14].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[15].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[16].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[17].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[19].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[18].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[21].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[22].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[23].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[24].acv_ac_ldc|adc_clk_cps ;
wire \address_gen[20].acv_ac_ldc|adc_clk_cps ;
wire \clock_gen[0].umem_ck_pad|auto_generated|dataout[0] ;
wire \mem_ck_source[0] ;
wire \clock_gen[0].leveled_dqs_clocks[0] ;
wire \clock_gen[0].leveled_dqs_clocks[1] ;
wire \clock_gen[0].leveled_dqs_clocks[2] ;
wire \clock_gen[0].leveled_dqs_clocks[3] ;

wire [3:0] \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ;

assign \clock_gen[0].leveled_dqs_clocks[0]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [0];
assign \clock_gen[0].leveled_dqs_clocks[1]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [1];
assign \clock_gen[0].leveled_dqs_clocks[2]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [2];
assign \clock_gen[0].leveled_dqs_clocks[3]  = \clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus [3];

terminal_qsys_hps_sdram_p0_acv_ldc \address_gen[0].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[0].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_23 \address_gen[8].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[8].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_22 \address_gen[7].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[7].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_21 \address_gen[6].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[6].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_20 \address_gen[5].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[5].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_19 \address_gen[4].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[4].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_18 \address_gen[3].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[3].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_17 \address_gen[2].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[2].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_11 \address_gen[1].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[1].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_6 \address_gen[15].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[15].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_5 \address_gen[14].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[14].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_4 \address_gen[13].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[13].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_3 \address_gen[12].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[12].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_2 \address_gen[11].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[11].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_1 \address_gen[10].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[10].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_24 \address_gen[9].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[9].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_15 \address_gen[23].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[23].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_14 \address_gen[22].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[22].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_13 \address_gen[21].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[21].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_12 \address_gen[20].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[20].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_10 \address_gen[19].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[19].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_9 \address_gen[18].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[18].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_8 \address_gen[17].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[17].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_7 \address_gen[16].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[16].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

terminal_qsys_hps_sdram_p0_clock_pair_generator \clock_gen[0].uclk_generator (
	.wire_pseudo_diffa_o_0(wire_pseudo_diffa_o_0),
	.wire_pseudo_diffa_obar_0(wire_pseudo_diffa_obar_0),
	.wire_pseudo_diffa_oeout_0(wire_pseudo_diffa_oeout_0),
	.wire_pseudo_diffa_oebout_0(wire_pseudo_diffa_oebout_0),
	.datain({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }));

terminal_qsys_altddio_out_1 \clock_gen[0].umem_ck_pad (
	.dataout({\clock_gen[0].umem_ck_pad|auto_generated|dataout[0] }),
	.datain_h({phy_ddio_ck_0}),
	.datain_l({phy_ddio_ck_1}),
	.outclock(\mem_ck_source[0] ));

terminal_qsys_hps_sdram_p0_generic_ddio_3 ureset_n_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk}),
	.dataout({dataout_unconnected_wire_14,dataout_unconnected_wire_13,dataout_unconnected_wire_12,dataout_unconnected_wire_11,dataout_unconnected_wire_10,dataout_unconnected_wire_9,dataout_unconnected_wire_8,dataout_unconnected_wire_7,dataout_unconnected_wire_6,
dataout_unconnected_wire_5,dataout_unconnected_wire_4,dataout_unconnected_wire_3,dataout_unconnected_wire_2,dataout_unconnected_wire_1,dataout_03}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[24].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_reset_n_3,phy_ddio_reset_n_2,phy_ddio_reset_n_1,phy_ddio_reset_n_0}));

terminal_qsys_hps_sdram_p0_generic_ddio_2 ucmd_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_1,dataout_unconnected_wire_13_1,dataout_unconnected_wire_12_1,dataout_unconnected_wire_11_1,dataout_unconnected_wire_10_1,dataout_unconnected_wire_9_1,dataout_unconnected_wire_8_1,dataout_unconnected_wire_7_1,
dataout_unconnected_wire_6_1,dataout_51,dataout_41,dataout_31,dataout_22,dataout_16,dataout_02}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[23].acv_ac_ldc|adc_clk_cps ,\address_gen[22].acv_ac_ldc|adc_clk_cps ,\address_gen[21].acv_ac_ldc|adc_clk_cps ,\address_gen[20].acv_ac_ldc|adc_clk_cps ,\address_gen[19].acv_ac_ldc|adc_clk_cps ,
\address_gen[18].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_we_n_3,phy_ddio_we_n_2,phy_ddio_we_n_1,phy_ddio_we_n_0,phy_ddio_cas_n_3,phy_ddio_cas_n_2,phy_ddio_cas_n_1,phy_ddio_cas_n_0,phy_ddio_ras_n_3,
phy_ddio_ras_n_2,phy_ddio_ras_n_1,phy_ddio_ras_n_0,phy_ddio_odt_3,phy_ddio_odt_2,phy_ddio_odt_1,phy_ddio_odt_0,phy_ddio_cke_3,phy_ddio_cke_2,phy_ddio_cke_1,phy_ddio_cke_0,phy_ddio_cs_n_3,phy_ddio_cs_n_2,phy_ddio_cs_n_1,phy_ddio_cs_n_0}));

terminal_qsys_hps_sdram_p0_generic_ddio_1 ubank_pad(
	.clk_hr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_unconnected_wire_14_2,dataout_unconnected_wire_13_2,dataout_unconnected_wire_12_2,dataout_unconnected_wire_11_2,dataout_unconnected_wire_10_2,dataout_unconnected_wire_9_2,dataout_unconnected_wire_8_2,dataout_unconnected_wire_7_2,
dataout_unconnected_wire_6_2,dataout_unconnected_wire_5_1,dataout_unconnected_wire_4_1,dataout_unconnected_wire_3_1,dataout_21,dataout_15,dataout_01}),
	.clk_fr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\address_gen[17].acv_ac_ldc|adc_clk_cps ,\address_gen[16].acv_ac_ldc|adc_clk_cps ,\address_gen[15].acv_ac_ldc|adc_clk_cps }),
	.datain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,phy_ddio_bank_11,phy_ddio_bank_10,phy_ddio_bank_9,phy_ddio_bank_8,phy_ddio_bank_7,phy_ddio_bank_6,phy_ddio_bank_5,
phy_ddio_bank_4,phy_ddio_bank_3,phy_ddio_bank_2,phy_ddio_bank_1,phy_ddio_bank_0}));

terminal_qsys_hps_sdram_p0_generic_ddio uaddress_pad(
	.clk_hr({afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk,afi_clk}),
	.dataout({dataout_14,dataout_13,dataout_12,dataout_11,dataout_10,dataout_9,dataout_8,dataout_7,dataout_6,dataout_5,dataout_4,dataout_3,dataout_2,dataout_1,dataout_0}),
	.clk_fr({\address_gen[14].acv_ac_ldc|adc_clk_cps ,\address_gen[13].acv_ac_ldc|adc_clk_cps ,\address_gen[12].acv_ac_ldc|adc_clk_cps ,\address_gen[11].acv_ac_ldc|adc_clk_cps ,\address_gen[10].acv_ac_ldc|adc_clk_cps ,\address_gen[9].acv_ac_ldc|adc_clk_cps ,
\address_gen[8].acv_ac_ldc|adc_clk_cps ,\address_gen[7].acv_ac_ldc|adc_clk_cps ,\address_gen[6].acv_ac_ldc|adc_clk_cps ,\address_gen[5].acv_ac_ldc|adc_clk_cps ,\address_gen[4].acv_ac_ldc|adc_clk_cps ,\address_gen[3].acv_ac_ldc|adc_clk_cps ,
\address_gen[2].acv_ac_ldc|adc_clk_cps ,\address_gen[1].acv_ac_ldc|adc_clk_cps ,\address_gen[0].acv_ac_ldc|adc_clk_cps }),
	.datain({phy_ddio_address_59,phy_ddio_address_58,phy_ddio_address_57,phy_ddio_address_56,phy_ddio_address_55,phy_ddio_address_54,phy_ddio_address_53,phy_ddio_address_52,phy_ddio_address_51,phy_ddio_address_50,phy_ddio_address_49,phy_ddio_address_48,phy_ddio_address_47,
phy_ddio_address_46,phy_ddio_address_45,phy_ddio_address_44,phy_ddio_address_43,phy_ddio_address_42,phy_ddio_address_41,phy_ddio_address_40,phy_ddio_address_39,phy_ddio_address_38,phy_ddio_address_37,phy_ddio_address_36,phy_ddio_address_35,phy_ddio_address_34,
phy_ddio_address_33,phy_ddio_address_32,phy_ddio_address_31,phy_ddio_address_30,phy_ddio_address_29,phy_ddio_address_28,phy_ddio_address_27,phy_ddio_address_26,phy_ddio_address_25,phy_ddio_address_24,phy_ddio_address_23,phy_ddio_address_22,phy_ddio_address_21,
phy_ddio_address_20,phy_ddio_address_19,phy_ddio_address_18,phy_ddio_address_17,phy_ddio_address_16,phy_ddio_address_15,phy_ddio_address_14,phy_ddio_address_13,phy_ddio_address_12,phy_ddio_address_11,phy_ddio_address_10,phy_ddio_address_9,phy_ddio_address_8,
phy_ddio_address_7,phy_ddio_address_6,phy_ddio_address_5,phy_ddio_address_4,phy_ddio_address_3,phy_ddio_address_2,phy_ddio_address_1,phy_ddio_address_0}));

terminal_qsys_hps_sdram_p0_acv_ldc_16 \address_gen[24].acv_ac_ldc (
	.pll_dqs_clk(afi_clk),
	.adc_clk_cps(\address_gen[24].acv_ac_ldc|adc_clk_cps ),
	.dll_phy_delayctrl({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}));

cyclonev_clk_phase_select \clock_gen[0].clk_phase_select_dqs (
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\clock_gen[0].leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(\mem_ck_source[0] ));
defparam \clock_gen[0].clk_phase_select_dqs .invert_phase = "false";
defparam \clock_gen[0].clk_phase_select_dqs .phase_setting = 0;
defparam \clock_gen[0].clk_phase_select_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].clk_phase_select_dqs .use_dqs_input = "false";
defparam \clock_gen[0].clk_phase_select_dqs .use_phasectrlin = "false";

cyclonev_leveling_delay_chain \clock_gen[0].leveling_delay_chain_dqs (
	.clkin(afi_clk),
	.delayctrlin({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.clkout(\clock_gen[0].leveling_delay_chain_dqs_CLKOUT_bus ));
defparam \clock_gen[0].leveling_delay_chain_dqs .physical_clock_source = "dqs";
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_delay_increment = 10;
defparam \clock_gen[0].leveling_delay_chain_dqs .sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_altddio_out_1 (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
inout 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_ddio_out_uqe auto_generated(
	.dataout({dataout[0]}),
	.datain_h({datain_h[0]}),
	.datain_l({datain_l[0]}),
	.outclock(outclock));

endmodule

module terminal_qsys_ddio_out_uqe (
	dataout,
	datain_h,
	datain_l,
	outclock)/* synthesis synthesis_greybox=0 */;
output 	[0:0] dataout;
input 	[0:0] datain_h;
input 	[0:0] datain_l;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "none";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_1 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_2 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_3 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_4 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_5 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_6 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_7 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_8 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_9 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_10 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_11 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_12 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_13 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_14 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_15 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_16 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_17 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_18 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_19 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_20 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_21 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_22 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_23 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_24 (
	pll_dqs_clk,
	adc_clk_cps,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
output 	adc_clk_cps;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_clk_phase_select clk_phase_select_addr_cmd(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(adc_clk_cps));
defparam clk_phase_select_addr_cmd.invert_phase = "true";
defparam clk_phase_select_addr_cmd.phase_setting = 0;
defparam clk_phase_select_addr_cmd.physical_clock_source = "add_cmd";
defparam clk_phase_select_addr_cmd.use_dqs_input = "false";
defparam clk_phase_select_addr_cmd.use_phasectrlin = "false";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_p0_clock_pair_generator (
	wire_pseudo_diffa_o_0,
	wire_pseudo_diffa_obar_0,
	wire_pseudo_diffa_oeout_0,
	wire_pseudo_diffa_oebout_0,
	datain)/* synthesis synthesis_greybox=0 */;
output 	wire_pseudo_diffa_o_0;
output 	wire_pseudo_diffa_obar_0;
output 	wire_pseudo_diffa_oeout_0;
output 	wire_pseudo_diffa_oebout_0;
input 	[0:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(datain[0]),
	.oein(gnd),
	.dtcin(gnd),
	.o(wire_pseudo_diffa_o_0),
	.obar(wire_pseudo_diffa_obar_0),
	.oeout(wire_pseudo_diffa_oeout_0),
	.oebout(wire_pseudo_diffa_oebout_0),
	.dtc(),
	.dtcbar());

endmodule

module terminal_qsys_hps_sdram_p0_generic_ddio (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[6].fr_data_lo ;
wire \acblock[6].fr_data_hi ;
wire \acblock[7].fr_data_lo ;
wire \acblock[7].fr_data_hi ;
wire \acblock[8].fr_data_lo ;
wire \acblock[8].fr_data_hi ;
wire \acblock[9].fr_data_lo ;
wire \acblock[9].fr_data_hi ;
wire \acblock[10].fr_data_lo ;
wire \acblock[10].fr_data_hi ;
wire \acblock[11].fr_data_lo ;
wire \acblock[11].fr_data_hi ;
wire \acblock[12].fr_data_lo ;
wire \acblock[12].fr_data_hi ;
wire \acblock[13].fr_data_lo ;
wire \acblock[13].fr_data_hi ;
wire \acblock[14].fr_data_lo ;
wire \acblock[14].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].ddio_out (
	.datainlo(\acblock[6].fr_data_lo ),
	.datainhi(\acblock[6].fr_data_hi ),
	.clkhi(clk_fr[6]),
	.clklo(clk_fr[6]),
	.muxsel(clk_fr[6]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[6]),
	.dfflo(),
	.dffhi());
defparam \acblock[6].ddio_out .async_mode = "none";
defparam \acblock[6].ddio_out .half_rate_mode = "false";
defparam \acblock[6].ddio_out .power_up = "low";
defparam \acblock[6].ddio_out .sync_mode = "none";
defparam \acblock[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].ddio_out (
	.datainlo(\acblock[7].fr_data_lo ),
	.datainhi(\acblock[7].fr_data_hi ),
	.clkhi(clk_fr[7]),
	.clklo(clk_fr[7]),
	.muxsel(clk_fr[7]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[7]),
	.dfflo(),
	.dffhi());
defparam \acblock[7].ddio_out .async_mode = "none";
defparam \acblock[7].ddio_out .half_rate_mode = "false";
defparam \acblock[7].ddio_out .power_up = "low";
defparam \acblock[7].ddio_out .sync_mode = "none";
defparam \acblock[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].ddio_out (
	.datainlo(\acblock[8].fr_data_lo ),
	.datainhi(\acblock[8].fr_data_hi ),
	.clkhi(clk_fr[8]),
	.clklo(clk_fr[8]),
	.muxsel(clk_fr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[8]),
	.dfflo(),
	.dffhi());
defparam \acblock[8].ddio_out .async_mode = "none";
defparam \acblock[8].ddio_out .half_rate_mode = "false";
defparam \acblock[8].ddio_out .power_up = "low";
defparam \acblock[8].ddio_out .sync_mode = "none";
defparam \acblock[8].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].ddio_out (
	.datainlo(\acblock[9].fr_data_lo ),
	.datainhi(\acblock[9].fr_data_hi ),
	.clkhi(clk_fr[9]),
	.clklo(clk_fr[9]),
	.muxsel(clk_fr[9]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[9]),
	.dfflo(),
	.dffhi());
defparam \acblock[9].ddio_out .async_mode = "none";
defparam \acblock[9].ddio_out .half_rate_mode = "false";
defparam \acblock[9].ddio_out .power_up = "low";
defparam \acblock[9].ddio_out .sync_mode = "none";
defparam \acblock[9].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].ddio_out (
	.datainlo(\acblock[10].fr_data_lo ),
	.datainhi(\acblock[10].fr_data_hi ),
	.clkhi(clk_fr[10]),
	.clklo(clk_fr[10]),
	.muxsel(clk_fr[10]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[10]),
	.dfflo(),
	.dffhi());
defparam \acblock[10].ddio_out .async_mode = "none";
defparam \acblock[10].ddio_out .half_rate_mode = "false";
defparam \acblock[10].ddio_out .power_up = "low";
defparam \acblock[10].ddio_out .sync_mode = "none";
defparam \acblock[10].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].ddio_out (
	.datainlo(\acblock[11].fr_data_lo ),
	.datainhi(\acblock[11].fr_data_hi ),
	.clkhi(clk_fr[11]),
	.clklo(clk_fr[11]),
	.muxsel(clk_fr[11]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[11]),
	.dfflo(),
	.dffhi());
defparam \acblock[11].ddio_out .async_mode = "none";
defparam \acblock[11].ddio_out .half_rate_mode = "false";
defparam \acblock[11].ddio_out .power_up = "low";
defparam \acblock[11].ddio_out .sync_mode = "none";
defparam \acblock[11].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].ddio_out (
	.datainlo(\acblock[12].fr_data_lo ),
	.datainhi(\acblock[12].fr_data_hi ),
	.clkhi(clk_fr[12]),
	.clklo(clk_fr[12]),
	.muxsel(clk_fr[12]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[12]),
	.dfflo(),
	.dffhi());
defparam \acblock[12].ddio_out .async_mode = "none";
defparam \acblock[12].ddio_out .half_rate_mode = "false";
defparam \acblock[12].ddio_out .power_up = "low";
defparam \acblock[12].ddio_out .sync_mode = "none";
defparam \acblock[12].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].ddio_out (
	.datainlo(\acblock[13].fr_data_lo ),
	.datainhi(\acblock[13].fr_data_hi ),
	.clkhi(clk_fr[13]),
	.clklo(clk_fr[13]),
	.muxsel(clk_fr[13]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[13]),
	.dfflo(),
	.dffhi());
defparam \acblock[13].ddio_out .async_mode = "none";
defparam \acblock[13].ddio_out .half_rate_mode = "false";
defparam \acblock[13].ddio_out .power_up = "low";
defparam \acblock[13].ddio_out .sync_mode = "none";
defparam \acblock[13].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].ddio_out (
	.datainlo(\acblock[14].fr_data_lo ),
	.datainhi(\acblock[14].fr_data_hi ),
	.clkhi(clk_fr[14]),
	.clklo(clk_fr[14]),
	.muxsel(clk_fr[14]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[14]),
	.dfflo(),
	.dffhi());
defparam \acblock[14].ddio_out .async_mode = "none";
defparam \acblock[14].ddio_out .half_rate_mode = "false";
defparam \acblock[14].ddio_out .power_up = "low";
defparam \acblock[14].ddio_out .sync_mode = "none";
defparam \acblock[14].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_lo (
	.datainlo(datain[27]),
	.datainhi(datain[25]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_lo .async_mode = "none";
defparam \acblock[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_lo .power_up = "low";
defparam \acblock[6].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[6].hr_to_fr_hi (
	.datainlo(datain[26]),
	.datainhi(datain[24]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[6].hr_to_fr_hi .async_mode = "none";
defparam \acblock[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[6].hr_to_fr_hi .power_up = "low";
defparam \acblock[6].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_lo (
	.datainlo(datain[31]),
	.datainhi(datain[29]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_lo .async_mode = "none";
defparam \acblock[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_lo .power_up = "low";
defparam \acblock[7].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[7].hr_to_fr_hi (
	.datainlo(datain[30]),
	.datainhi(datain[28]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[7].hr_to_fr_hi .async_mode = "none";
defparam \acblock[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[7].hr_to_fr_hi .power_up = "low";
defparam \acblock[7].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_lo (
	.datainlo(datain[35]),
	.datainhi(datain[33]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_lo .async_mode = "none";
defparam \acblock[8].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_lo .power_up = "low";
defparam \acblock[8].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[8].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[8].hr_to_fr_hi (
	.datainlo(datain[34]),
	.datainhi(datain[32]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[8].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[8].hr_to_fr_hi .async_mode = "none";
defparam \acblock[8].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[8].hr_to_fr_hi .power_up = "low";
defparam \acblock[8].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[8].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_lo (
	.datainlo(datain[39]),
	.datainhi(datain[37]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_lo .async_mode = "none";
defparam \acblock[9].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_lo .power_up = "low";
defparam \acblock[9].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[9].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[9].hr_to_fr_hi (
	.datainlo(datain[38]),
	.datainhi(datain[36]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[9].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[9].hr_to_fr_hi .async_mode = "none";
defparam \acblock[9].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[9].hr_to_fr_hi .power_up = "low";
defparam \acblock[9].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[9].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_lo (
	.datainlo(datain[43]),
	.datainhi(datain[41]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_lo .async_mode = "none";
defparam \acblock[10].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_lo .power_up = "low";
defparam \acblock[10].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[10].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[10].hr_to_fr_hi (
	.datainlo(datain[42]),
	.datainhi(datain[40]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[10].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[10].hr_to_fr_hi .async_mode = "none";
defparam \acblock[10].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[10].hr_to_fr_hi .power_up = "low";
defparam \acblock[10].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[10].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_lo (
	.datainlo(datain[47]),
	.datainhi(datain[45]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_lo .async_mode = "none";
defparam \acblock[11].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_lo .power_up = "low";
defparam \acblock[11].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[11].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[11].hr_to_fr_hi (
	.datainlo(datain[46]),
	.datainhi(datain[44]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[11].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[11].hr_to_fr_hi .async_mode = "none";
defparam \acblock[11].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[11].hr_to_fr_hi .power_up = "low";
defparam \acblock[11].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[11].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_lo (
	.datainlo(datain[51]),
	.datainhi(datain[49]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_lo .async_mode = "none";
defparam \acblock[12].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_lo .power_up = "low";
defparam \acblock[12].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[12].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[12].hr_to_fr_hi (
	.datainlo(datain[50]),
	.datainhi(datain[48]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[12].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[12].hr_to_fr_hi .async_mode = "none";
defparam \acblock[12].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[12].hr_to_fr_hi .power_up = "low";
defparam \acblock[12].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[12].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_lo (
	.datainlo(datain[55]),
	.datainhi(datain[53]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_lo .async_mode = "none";
defparam \acblock[13].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_lo .power_up = "low";
defparam \acblock[13].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[13].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[13].hr_to_fr_hi (
	.datainlo(datain[54]),
	.datainhi(datain[52]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[13].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[13].hr_to_fr_hi .async_mode = "none";
defparam \acblock[13].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[13].hr_to_fr_hi .power_up = "low";
defparam \acblock[13].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[13].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_lo (
	.datainlo(datain[59]),
	.datainhi(datain[57]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_lo .async_mode = "none";
defparam \acblock[14].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_lo .power_up = "low";
defparam \acblock[14].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[14].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[14].hr_to_fr_hi (
	.datainlo(datain[58]),
	.datainhi(datain[56]),
	.clkhi(clk_hr[8]),
	.clklo(clk_hr[8]),
	.muxsel(clk_hr[8]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[14].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[14].hr_to_fr_hi .async_mode = "none";
defparam \acblock[14].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[14].hr_to_fr_hi .power_up = "low";
defparam \acblock[14].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[14].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_generic_ddio_1 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_generic_ddio_2 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[1].fr_data_lo ;
wire \acblock[1].fr_data_hi ;
wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;
wire \acblock[3].fr_data_lo ;
wire \acblock[3].fr_data_hi ;
wire \acblock[4].fr_data_lo ;
wire \acblock[4].fr_data_hi ;
wire \acblock[5].fr_data_lo ;
wire \acblock[5].fr_data_hi ;
wire \acblock[2].fr_data_lo ;
wire \acblock[2].fr_data_hi ;


cyclonev_ddio_out \acblock[1].ddio_out (
	.datainlo(\acblock[1].fr_data_lo ),
	.datainhi(\acblock[1].fr_data_hi ),
	.clkhi(clk_fr[1]),
	.clklo(clk_fr[1]),
	.muxsel(clk_fr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \acblock[1].ddio_out .async_mode = "none";
defparam \acblock[1].ddio_out .half_rate_mode = "false";
defparam \acblock[1].ddio_out .power_up = "low";
defparam \acblock[1].ddio_out .sync_mode = "none";
defparam \acblock[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].ddio_out (
	.datainlo(\acblock[3].fr_data_lo ),
	.datainhi(\acblock[3].fr_data_hi ),
	.clkhi(clk_fr[3]),
	.clklo(clk_fr[3]),
	.muxsel(clk_fr[3]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \acblock[3].ddio_out .async_mode = "none";
defparam \acblock[3].ddio_out .half_rate_mode = "false";
defparam \acblock[3].ddio_out .power_up = "low";
defparam \acblock[3].ddio_out .sync_mode = "none";
defparam \acblock[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].ddio_out (
	.datainlo(\acblock[4].fr_data_lo ),
	.datainhi(\acblock[4].fr_data_hi ),
	.clkhi(clk_fr[4]),
	.clklo(clk_fr[4]),
	.muxsel(clk_fr[4]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[4]),
	.dfflo(),
	.dffhi());
defparam \acblock[4].ddio_out .async_mode = "none";
defparam \acblock[4].ddio_out .half_rate_mode = "false";
defparam \acblock[4].ddio_out .power_up = "low";
defparam \acblock[4].ddio_out .sync_mode = "none";
defparam \acblock[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].ddio_out (
	.datainlo(\acblock[5].fr_data_lo ),
	.datainhi(\acblock[5].fr_data_hi ),
	.clkhi(clk_fr[5]),
	.clklo(clk_fr[5]),
	.muxsel(clk_fr[5]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[5]),
	.dfflo(),
	.dffhi());
defparam \acblock[5].ddio_out .async_mode = "none";
defparam \acblock[5].ddio_out .half_rate_mode = "false";
defparam \acblock[5].ddio_out .power_up = "low";
defparam \acblock[5].ddio_out .sync_mode = "none";
defparam \acblock[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].ddio_out (
	.datainlo(\acblock[2].fr_data_lo ),
	.datainhi(\acblock[2].fr_data_hi ),
	.clkhi(clk_fr[2]),
	.clklo(clk_fr[2]),
	.muxsel(clk_fr[2]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \acblock[2].ddio_out .async_mode = "none";
defparam \acblock[2].ddio_out .half_rate_mode = "false";
defparam \acblock[2].ddio_out .power_up = "low";
defparam \acblock[2].ddio_out .sync_mode = "none";
defparam \acblock[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_lo (
	.datainlo(datain[7]),
	.datainhi(datain[5]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_lo .async_mode = "none";
defparam \acblock[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_lo .power_up = "low";
defparam \acblock[1].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[1].hr_to_fr_hi (
	.datainlo(datain[6]),
	.datainhi(datain[4]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[1].hr_to_fr_hi .async_mode = "none";
defparam \acblock[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[1].hr_to_fr_hi .power_up = "low";
defparam \acblock[1].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_lo (
	.datainlo(datain[15]),
	.datainhi(datain[13]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_lo .async_mode = "none";
defparam \acblock[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_lo .power_up = "low";
defparam \acblock[3].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[3].hr_to_fr_hi (
	.datainlo(datain[14]),
	.datainhi(datain[12]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[3].hr_to_fr_hi .async_mode = "none";
defparam \acblock[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[3].hr_to_fr_hi .power_up = "low";
defparam \acblock[3].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_lo (
	.datainlo(datain[19]),
	.datainhi(datain[17]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_lo .async_mode = "none";
defparam \acblock[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_lo .power_up = "low";
defparam \acblock[4].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[4].hr_to_fr_hi (
	.datainlo(datain[18]),
	.datainhi(datain[16]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[4].hr_to_fr_hi .async_mode = "none";
defparam \acblock[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[4].hr_to_fr_hi .power_up = "low";
defparam \acblock[4].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_lo (
	.datainlo(datain[23]),
	.datainhi(datain[21]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_lo .async_mode = "none";
defparam \acblock[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_lo .power_up = "low";
defparam \acblock[5].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[5].hr_to_fr_hi (
	.datainlo(datain[22]),
	.datainhi(datain[20]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[5].hr_to_fr_hi .async_mode = "none";
defparam \acblock[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[5].hr_to_fr_hi .power_up = "low";
defparam \acblock[5].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_lo (
	.datainlo(datain[11]),
	.datainhi(datain[9]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_lo .async_mode = "none";
defparam \acblock[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_lo .power_up = "low";
defparam \acblock[2].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[2].hr_to_fr_hi (
	.datainlo(datain[10]),
	.datainhi(datain[8]),
	.clkhi(clk_hr[1]),
	.clklo(clk_hr[1]),
	.muxsel(clk_hr[1]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[2].hr_to_fr_hi .async_mode = "none";
defparam \acblock[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[2].hr_to_fr_hi .power_up = "low";
defparam \acblock[2].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[2].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_generic_ddio_3 (
	clk_hr,
	dataout,
	clk_fr,
	datain)/* synthesis synthesis_greybox=0 */;
input 	[14:0] clk_hr;
output 	[14:0] dataout;
input 	[14:0] clk_fr;
input 	[59:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \acblock[0].fr_data_lo ;
wire \acblock[0].fr_data_hi ;


cyclonev_ddio_out \acblock[0].ddio_out (
	.datainlo(\acblock[0].fr_data_lo ),
	.datainhi(\acblock[0].fr_data_hi ),
	.clkhi(clk_fr[0]),
	.clklo(clk_fr[0]),
	.muxsel(clk_fr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \acblock[0].ddio_out .async_mode = "none";
defparam \acblock[0].ddio_out .half_rate_mode = "false";
defparam \acblock[0].ddio_out .power_up = "low";
defparam \acblock[0].ddio_out .sync_mode = "none";
defparam \acblock[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_lo (
	.datainlo(datain[3]),
	.datainhi(datain[1]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_lo .async_mode = "none";
defparam \acblock[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_lo .power_up = "low";
defparam \acblock[0].hr_to_fr_lo .sync_mode = "none";
defparam \acblock[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \acblock[0].hr_to_fr_hi (
	.datainlo(datain[2]),
	.datainhi(datain[0]),
	.clkhi(clk_hr[0]),
	.clklo(clk_hr[0]),
	.muxsel(clk_hr[0]),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(\acblock[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \acblock[0].hr_to_fr_hi .async_mode = "none";
defparam \acblock[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \acblock[0].hr_to_fr_hi .power_up = "low";
defparam \acblock[0].hr_to_fr_hi .sync_mode = "none";
defparam \acblock[0].hr_to_fr_hi .use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_altdqdqs (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_0,
	phy_ddio_dmdout_1,
	phy_ddio_dmdout_2,
	phy_ddio_dmdout_3,
	phy_ddio_dqdout_0,
	phy_ddio_dqdout_1,
	phy_ddio_dqdout_2,
	phy_ddio_dqdout_3,
	phy_ddio_dqdout_4,
	phy_ddio_dqdout_5,
	phy_ddio_dqdout_6,
	phy_ddio_dqdout_7,
	phy_ddio_dqdout_8,
	phy_ddio_dqdout_9,
	phy_ddio_dqdout_10,
	phy_ddio_dqdout_11,
	phy_ddio_dqdout_12,
	phy_ddio_dqdout_13,
	phy_ddio_dqdout_14,
	phy_ddio_dqdout_15,
	phy_ddio_dqdout_16,
	phy_ddio_dqdout_17,
	phy_ddio_dqdout_18,
	phy_ddio_dqdout_19,
	phy_ddio_dqdout_20,
	phy_ddio_dqdout_21,
	phy_ddio_dqdout_22,
	phy_ddio_dqdout_23,
	phy_ddio_dqdout_24,
	phy_ddio_dqdout_25,
	phy_ddio_dqdout_26,
	phy_ddio_dqdout_27,
	phy_ddio_dqdout_28,
	phy_ddio_dqdout_29,
	phy_ddio_dqdout_30,
	phy_ddio_dqdout_31,
	phy_ddio_dqoe_0,
	phy_ddio_dqoe_1,
	phy_ddio_dqoe_2,
	phy_ddio_dqoe_3,
	phy_ddio_dqoe_4,
	phy_ddio_dqoe_5,
	phy_ddio_dqoe_6,
	phy_ddio_dqoe_7,
	phy_ddio_dqoe_8,
	phy_ddio_dqoe_9,
	phy_ddio_dqoe_10,
	phy_ddio_dqoe_11,
	phy_ddio_dqoe_12,
	phy_ddio_dqoe_13,
	phy_ddio_dqoe_14,
	phy_ddio_dqoe_15,
	phy_ddio_dqs_dout_0,
	phy_ddio_dqs_dout_1,
	phy_ddio_dqs_dout_2,
	phy_ddio_dqs_dout_3,
	phy_ddio_dqslogic_aclr_fifoctrl_0,
	phy_ddio_dqslogic_aclr_pstamble_0,
	phy_ddio_dqslogic_dqsena_0,
	phy_ddio_dqslogic_dqsena_1,
	phy_ddio_dqslogic_fiforeset_0,
	phy_ddio_dqslogic_incrdataen_0,
	phy_ddio_dqslogic_incrdataen_1,
	phy_ddio_dqslogic_incwrptr_0,
	phy_ddio_dqslogic_incwrptr_1,
	phy_ddio_dqslogic_oct_0,
	phy_ddio_dqslogic_oct_1,
	phy_ddio_dqslogic_readlatency_0,
	phy_ddio_dqslogic_readlatency_1,
	phy_ddio_dqslogic_readlatency_2,
	phy_ddio_dqslogic_readlatency_3,
	phy_ddio_dqslogic_readlatency_4,
	phy_ddio_dqs_oe_0,
	phy_ddio_dqs_oe_1,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_0;
input 	phy_ddio_dmdout_1;
input 	phy_ddio_dmdout_2;
input 	phy_ddio_dmdout_3;
input 	phy_ddio_dqdout_0;
input 	phy_ddio_dqdout_1;
input 	phy_ddio_dqdout_2;
input 	phy_ddio_dqdout_3;
input 	phy_ddio_dqdout_4;
input 	phy_ddio_dqdout_5;
input 	phy_ddio_dqdout_6;
input 	phy_ddio_dqdout_7;
input 	phy_ddio_dqdout_8;
input 	phy_ddio_dqdout_9;
input 	phy_ddio_dqdout_10;
input 	phy_ddio_dqdout_11;
input 	phy_ddio_dqdout_12;
input 	phy_ddio_dqdout_13;
input 	phy_ddio_dqdout_14;
input 	phy_ddio_dqdout_15;
input 	phy_ddio_dqdout_16;
input 	phy_ddio_dqdout_17;
input 	phy_ddio_dqdout_18;
input 	phy_ddio_dqdout_19;
input 	phy_ddio_dqdout_20;
input 	phy_ddio_dqdout_21;
input 	phy_ddio_dqdout_22;
input 	phy_ddio_dqdout_23;
input 	phy_ddio_dqdout_24;
input 	phy_ddio_dqdout_25;
input 	phy_ddio_dqdout_26;
input 	phy_ddio_dqdout_27;
input 	phy_ddio_dqdout_28;
input 	phy_ddio_dqdout_29;
input 	phy_ddio_dqdout_30;
input 	phy_ddio_dqdout_31;
input 	phy_ddio_dqoe_0;
input 	phy_ddio_dqoe_1;
input 	phy_ddio_dqoe_2;
input 	phy_ddio_dqoe_3;
input 	phy_ddio_dqoe_4;
input 	phy_ddio_dqoe_5;
input 	phy_ddio_dqoe_6;
input 	phy_ddio_dqoe_7;
input 	phy_ddio_dqoe_8;
input 	phy_ddio_dqoe_9;
input 	phy_ddio_dqoe_10;
input 	phy_ddio_dqoe_11;
input 	phy_ddio_dqoe_12;
input 	phy_ddio_dqoe_13;
input 	phy_ddio_dqoe_14;
input 	phy_ddio_dqoe_15;
input 	phy_ddio_dqs_dout_0;
input 	phy_ddio_dqs_dout_1;
input 	phy_ddio_dqs_dout_2;
input 	phy_ddio_dqs_dout_3;
input 	phy_ddio_dqslogic_aclr_fifoctrl_0;
input 	phy_ddio_dqslogic_aclr_pstamble_0;
input 	phy_ddio_dqslogic_dqsena_0;
input 	phy_ddio_dqslogic_dqsena_1;
input 	phy_ddio_dqslogic_fiforeset_0;
input 	phy_ddio_dqslogic_incrdataen_0;
input 	phy_ddio_dqslogic_incrdataen_1;
input 	phy_ddio_dqslogic_incwrptr_0;
input 	phy_ddio_dqslogic_incwrptr_1;
input 	phy_ddio_dqslogic_oct_0;
input 	phy_ddio_dqslogic_oct_1;
input 	phy_ddio_dqslogic_readlatency_0;
input 	phy_ddio_dqslogic_readlatency_1;
input 	phy_ddio_dqslogic_readlatency_2;
input 	phy_ddio_dqslogic_readlatency_3;
input 	phy_ddio_dqslogic_readlatency_4;
input 	phy_ddio_dqs_oe_0;
input 	phy_ddio_dqs_oe_1;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_3,phy_ddio_dmdout_2,phy_ddio_dmdout_1,phy_ddio_dmdout_0}),
	.write_data_in({phy_ddio_dqdout_31,phy_ddio_dqdout_30,phy_ddio_dqdout_29,phy_ddio_dqdout_28,phy_ddio_dqdout_27,phy_ddio_dqdout_26,phy_ddio_dqdout_25,phy_ddio_dqdout_24,phy_ddio_dqdout_23,phy_ddio_dqdout_22,phy_ddio_dqdout_21,phy_ddio_dqdout_20,phy_ddio_dqdout_19,phy_ddio_dqdout_18,
phy_ddio_dqdout_17,phy_ddio_dqdout_16,phy_ddio_dqdout_15,phy_ddio_dqdout_14,phy_ddio_dqdout_13,phy_ddio_dqdout_12,phy_ddio_dqdout_11,phy_ddio_dqdout_10,phy_ddio_dqdout_9,phy_ddio_dqdout_8,phy_ddio_dqdout_7,phy_ddio_dqdout_6,phy_ddio_dqdout_5,phy_ddio_dqdout_4,
phy_ddio_dqdout_3,phy_ddio_dqdout_2,phy_ddio_dqdout_1,phy_ddio_dqdout_0}),
	.write_oe_in({phy_ddio_dqoe_15,phy_ddio_dqoe_14,phy_ddio_dqoe_13,phy_ddio_dqoe_12,phy_ddio_dqoe_11,phy_ddio_dqoe_10,phy_ddio_dqoe_9,phy_ddio_dqoe_8,phy_ddio_dqoe_7,phy_ddio_dqoe_6,phy_ddio_dqoe_5,phy_ddio_dqoe_4,phy_ddio_dqoe_3,phy_ddio_dqoe_2,phy_ddio_dqoe_1,phy_ddio_dqoe_0}),
	.write_strobe({phy_ddio_dqs_dout_3,phy_ddio_dqs_dout_2,phy_ddio_dqs_dout_1,phy_ddio_dqs_dout_0}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_0),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_0),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_1,phy_ddio_dqslogic_dqsena_0}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_0),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_1,phy_ddio_dqslogic_incrdataen_0}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_1,phy_ddio_dqslogic_incwrptr_0}),
	.oct_ena_in({phy_ddio_dqslogic_oct_1,phy_ddio_dqslogic_oct_0}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_4,phy_ddio_dqslogic_readlatency_3,phy_ddio_dqslogic_readlatency_2,phy_ddio_dqslogic_readlatency_1,phy_ddio_dqslogic_readlatency_0}),
	.output_strobe_ena({phy_ddio_dqs_oe_1,phy_ddio_dqs_oe_0}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_altdqdqs_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_4,
	phy_ddio_dmdout_5,
	phy_ddio_dmdout_6,
	phy_ddio_dmdout_7,
	phy_ddio_dqdout_36,
	phy_ddio_dqdout_37,
	phy_ddio_dqdout_38,
	phy_ddio_dqdout_39,
	phy_ddio_dqdout_40,
	phy_ddio_dqdout_41,
	phy_ddio_dqdout_42,
	phy_ddio_dqdout_43,
	phy_ddio_dqdout_44,
	phy_ddio_dqdout_45,
	phy_ddio_dqdout_46,
	phy_ddio_dqdout_47,
	phy_ddio_dqdout_48,
	phy_ddio_dqdout_49,
	phy_ddio_dqdout_50,
	phy_ddio_dqdout_51,
	phy_ddio_dqdout_52,
	phy_ddio_dqdout_53,
	phy_ddio_dqdout_54,
	phy_ddio_dqdout_55,
	phy_ddio_dqdout_56,
	phy_ddio_dqdout_57,
	phy_ddio_dqdout_58,
	phy_ddio_dqdout_59,
	phy_ddio_dqdout_60,
	phy_ddio_dqdout_61,
	phy_ddio_dqdout_62,
	phy_ddio_dqdout_63,
	phy_ddio_dqdout_64,
	phy_ddio_dqdout_65,
	phy_ddio_dqdout_66,
	phy_ddio_dqdout_67,
	phy_ddio_dqoe_18,
	phy_ddio_dqoe_19,
	phy_ddio_dqoe_20,
	phy_ddio_dqoe_21,
	phy_ddio_dqoe_22,
	phy_ddio_dqoe_23,
	phy_ddio_dqoe_24,
	phy_ddio_dqoe_25,
	phy_ddio_dqoe_26,
	phy_ddio_dqoe_27,
	phy_ddio_dqoe_28,
	phy_ddio_dqoe_29,
	phy_ddio_dqoe_30,
	phy_ddio_dqoe_31,
	phy_ddio_dqoe_32,
	phy_ddio_dqoe_33,
	phy_ddio_dqs_dout_4,
	phy_ddio_dqs_dout_5,
	phy_ddio_dqs_dout_6,
	phy_ddio_dqs_dout_7,
	phy_ddio_dqslogic_aclr_fifoctrl_1,
	phy_ddio_dqslogic_aclr_pstamble_1,
	phy_ddio_dqslogic_dqsena_2,
	phy_ddio_dqslogic_dqsena_3,
	phy_ddio_dqslogic_fiforeset_1,
	phy_ddio_dqslogic_incrdataen_2,
	phy_ddio_dqslogic_incrdataen_3,
	phy_ddio_dqslogic_incwrptr_2,
	phy_ddio_dqslogic_incwrptr_3,
	phy_ddio_dqslogic_oct_2,
	phy_ddio_dqslogic_oct_3,
	phy_ddio_dqslogic_readlatency_5,
	phy_ddio_dqslogic_readlatency_6,
	phy_ddio_dqslogic_readlatency_7,
	phy_ddio_dqslogic_readlatency_8,
	phy_ddio_dqslogic_readlatency_9,
	phy_ddio_dqs_oe_2,
	phy_ddio_dqs_oe_3,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_4;
input 	phy_ddio_dmdout_5;
input 	phy_ddio_dmdout_6;
input 	phy_ddio_dmdout_7;
input 	phy_ddio_dqdout_36;
input 	phy_ddio_dqdout_37;
input 	phy_ddio_dqdout_38;
input 	phy_ddio_dqdout_39;
input 	phy_ddio_dqdout_40;
input 	phy_ddio_dqdout_41;
input 	phy_ddio_dqdout_42;
input 	phy_ddio_dqdout_43;
input 	phy_ddio_dqdout_44;
input 	phy_ddio_dqdout_45;
input 	phy_ddio_dqdout_46;
input 	phy_ddio_dqdout_47;
input 	phy_ddio_dqdout_48;
input 	phy_ddio_dqdout_49;
input 	phy_ddio_dqdout_50;
input 	phy_ddio_dqdout_51;
input 	phy_ddio_dqdout_52;
input 	phy_ddio_dqdout_53;
input 	phy_ddio_dqdout_54;
input 	phy_ddio_dqdout_55;
input 	phy_ddio_dqdout_56;
input 	phy_ddio_dqdout_57;
input 	phy_ddio_dqdout_58;
input 	phy_ddio_dqdout_59;
input 	phy_ddio_dqdout_60;
input 	phy_ddio_dqdout_61;
input 	phy_ddio_dqdout_62;
input 	phy_ddio_dqdout_63;
input 	phy_ddio_dqdout_64;
input 	phy_ddio_dqdout_65;
input 	phy_ddio_dqdout_66;
input 	phy_ddio_dqdout_67;
input 	phy_ddio_dqoe_18;
input 	phy_ddio_dqoe_19;
input 	phy_ddio_dqoe_20;
input 	phy_ddio_dqoe_21;
input 	phy_ddio_dqoe_22;
input 	phy_ddio_dqoe_23;
input 	phy_ddio_dqoe_24;
input 	phy_ddio_dqoe_25;
input 	phy_ddio_dqoe_26;
input 	phy_ddio_dqoe_27;
input 	phy_ddio_dqoe_28;
input 	phy_ddio_dqoe_29;
input 	phy_ddio_dqoe_30;
input 	phy_ddio_dqoe_31;
input 	phy_ddio_dqoe_32;
input 	phy_ddio_dqoe_33;
input 	phy_ddio_dqs_dout_4;
input 	phy_ddio_dqs_dout_5;
input 	phy_ddio_dqs_dout_6;
input 	phy_ddio_dqs_dout_7;
input 	phy_ddio_dqslogic_aclr_fifoctrl_1;
input 	phy_ddio_dqslogic_aclr_pstamble_1;
input 	phy_ddio_dqslogic_dqsena_2;
input 	phy_ddio_dqslogic_dqsena_3;
input 	phy_ddio_dqslogic_fiforeset_1;
input 	phy_ddio_dqslogic_incrdataen_2;
input 	phy_ddio_dqslogic_incrdataen_3;
input 	phy_ddio_dqslogic_incwrptr_2;
input 	phy_ddio_dqslogic_incwrptr_3;
input 	phy_ddio_dqslogic_oct_2;
input 	phy_ddio_dqslogic_oct_3;
input 	phy_ddio_dqslogic_readlatency_5;
input 	phy_ddio_dqslogic_readlatency_6;
input 	phy_ddio_dqslogic_readlatency_7;
input 	phy_ddio_dqslogic_readlatency_8;
input 	phy_ddio_dqslogic_readlatency_9;
input 	phy_ddio_dqs_oe_2;
input 	phy_ddio_dqs_oe_3;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_7,phy_ddio_dmdout_6,phy_ddio_dmdout_5,phy_ddio_dmdout_4}),
	.write_data_in({phy_ddio_dqdout_67,phy_ddio_dqdout_66,phy_ddio_dqdout_65,phy_ddio_dqdout_64,phy_ddio_dqdout_63,phy_ddio_dqdout_62,phy_ddio_dqdout_61,phy_ddio_dqdout_60,phy_ddio_dqdout_59,phy_ddio_dqdout_58,phy_ddio_dqdout_57,phy_ddio_dqdout_56,phy_ddio_dqdout_55,phy_ddio_dqdout_54,
phy_ddio_dqdout_53,phy_ddio_dqdout_52,phy_ddio_dqdout_51,phy_ddio_dqdout_50,phy_ddio_dqdout_49,phy_ddio_dqdout_48,phy_ddio_dqdout_47,phy_ddio_dqdout_46,phy_ddio_dqdout_45,phy_ddio_dqdout_44,phy_ddio_dqdout_43,phy_ddio_dqdout_42,phy_ddio_dqdout_41,phy_ddio_dqdout_40,
phy_ddio_dqdout_39,phy_ddio_dqdout_38,phy_ddio_dqdout_37,phy_ddio_dqdout_36}),
	.write_oe_in({phy_ddio_dqoe_33,phy_ddio_dqoe_32,phy_ddio_dqoe_31,phy_ddio_dqoe_30,phy_ddio_dqoe_29,phy_ddio_dqoe_28,phy_ddio_dqoe_27,phy_ddio_dqoe_26,phy_ddio_dqoe_25,phy_ddio_dqoe_24,phy_ddio_dqoe_23,phy_ddio_dqoe_22,phy_ddio_dqoe_21,phy_ddio_dqoe_20,phy_ddio_dqoe_19,phy_ddio_dqoe_18}),
	.write_strobe({phy_ddio_dqs_dout_7,phy_ddio_dqs_dout_6,phy_ddio_dqs_dout_5,phy_ddio_dqs_dout_4}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_1),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_1),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_3,phy_ddio_dqslogic_dqsena_2}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_1),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_3,phy_ddio_dqslogic_incrdataen_2}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_3,phy_ddio_dqslogic_incwrptr_2}),
	.oct_ena_in({phy_ddio_dqslogic_oct_3,phy_ddio_dqslogic_oct_2}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_9,phy_ddio_dqslogic_readlatency_8,phy_ddio_dqslogic_readlatency_7,phy_ddio_dqslogic_readlatency_6,phy_ddio_dqslogic_readlatency_5}),
	.output_strobe_ena({phy_ddio_dqs_oe_3,phy_ddio_dqs_oe_2}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_1 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_altdqdqs_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_8,
	phy_ddio_dmdout_9,
	phy_ddio_dmdout_10,
	phy_ddio_dmdout_11,
	phy_ddio_dqdout_72,
	phy_ddio_dqdout_73,
	phy_ddio_dqdout_74,
	phy_ddio_dqdout_75,
	phy_ddio_dqdout_76,
	phy_ddio_dqdout_77,
	phy_ddio_dqdout_78,
	phy_ddio_dqdout_79,
	phy_ddio_dqdout_80,
	phy_ddio_dqdout_81,
	phy_ddio_dqdout_82,
	phy_ddio_dqdout_83,
	phy_ddio_dqdout_84,
	phy_ddio_dqdout_85,
	phy_ddio_dqdout_86,
	phy_ddio_dqdout_87,
	phy_ddio_dqdout_88,
	phy_ddio_dqdout_89,
	phy_ddio_dqdout_90,
	phy_ddio_dqdout_91,
	phy_ddio_dqdout_92,
	phy_ddio_dqdout_93,
	phy_ddio_dqdout_94,
	phy_ddio_dqdout_95,
	phy_ddio_dqdout_96,
	phy_ddio_dqdout_97,
	phy_ddio_dqdout_98,
	phy_ddio_dqdout_99,
	phy_ddio_dqdout_100,
	phy_ddio_dqdout_101,
	phy_ddio_dqdout_102,
	phy_ddio_dqdout_103,
	phy_ddio_dqoe_36,
	phy_ddio_dqoe_37,
	phy_ddio_dqoe_38,
	phy_ddio_dqoe_39,
	phy_ddio_dqoe_40,
	phy_ddio_dqoe_41,
	phy_ddio_dqoe_42,
	phy_ddio_dqoe_43,
	phy_ddio_dqoe_44,
	phy_ddio_dqoe_45,
	phy_ddio_dqoe_46,
	phy_ddio_dqoe_47,
	phy_ddio_dqoe_48,
	phy_ddio_dqoe_49,
	phy_ddio_dqoe_50,
	phy_ddio_dqoe_51,
	phy_ddio_dqs_dout_8,
	phy_ddio_dqs_dout_9,
	phy_ddio_dqs_dout_10,
	phy_ddio_dqs_dout_11,
	phy_ddio_dqslogic_aclr_fifoctrl_2,
	phy_ddio_dqslogic_aclr_pstamble_2,
	phy_ddio_dqslogic_dqsena_4,
	phy_ddio_dqslogic_dqsena_5,
	phy_ddio_dqslogic_fiforeset_2,
	phy_ddio_dqslogic_incrdataen_4,
	phy_ddio_dqslogic_incrdataen_5,
	phy_ddio_dqslogic_incwrptr_4,
	phy_ddio_dqslogic_incwrptr_5,
	phy_ddio_dqslogic_oct_4,
	phy_ddio_dqslogic_oct_5,
	phy_ddio_dqslogic_readlatency_10,
	phy_ddio_dqslogic_readlatency_11,
	phy_ddio_dqslogic_readlatency_12,
	phy_ddio_dqslogic_readlatency_13,
	phy_ddio_dqslogic_readlatency_14,
	phy_ddio_dqs_oe_4,
	phy_ddio_dqs_oe_5,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_8;
input 	phy_ddio_dmdout_9;
input 	phy_ddio_dmdout_10;
input 	phy_ddio_dmdout_11;
input 	phy_ddio_dqdout_72;
input 	phy_ddio_dqdout_73;
input 	phy_ddio_dqdout_74;
input 	phy_ddio_dqdout_75;
input 	phy_ddio_dqdout_76;
input 	phy_ddio_dqdout_77;
input 	phy_ddio_dqdout_78;
input 	phy_ddio_dqdout_79;
input 	phy_ddio_dqdout_80;
input 	phy_ddio_dqdout_81;
input 	phy_ddio_dqdout_82;
input 	phy_ddio_dqdout_83;
input 	phy_ddio_dqdout_84;
input 	phy_ddio_dqdout_85;
input 	phy_ddio_dqdout_86;
input 	phy_ddio_dqdout_87;
input 	phy_ddio_dqdout_88;
input 	phy_ddio_dqdout_89;
input 	phy_ddio_dqdout_90;
input 	phy_ddio_dqdout_91;
input 	phy_ddio_dqdout_92;
input 	phy_ddio_dqdout_93;
input 	phy_ddio_dqdout_94;
input 	phy_ddio_dqdout_95;
input 	phy_ddio_dqdout_96;
input 	phy_ddio_dqdout_97;
input 	phy_ddio_dqdout_98;
input 	phy_ddio_dqdout_99;
input 	phy_ddio_dqdout_100;
input 	phy_ddio_dqdout_101;
input 	phy_ddio_dqdout_102;
input 	phy_ddio_dqdout_103;
input 	phy_ddio_dqoe_36;
input 	phy_ddio_dqoe_37;
input 	phy_ddio_dqoe_38;
input 	phy_ddio_dqoe_39;
input 	phy_ddio_dqoe_40;
input 	phy_ddio_dqoe_41;
input 	phy_ddio_dqoe_42;
input 	phy_ddio_dqoe_43;
input 	phy_ddio_dqoe_44;
input 	phy_ddio_dqoe_45;
input 	phy_ddio_dqoe_46;
input 	phy_ddio_dqoe_47;
input 	phy_ddio_dqoe_48;
input 	phy_ddio_dqoe_49;
input 	phy_ddio_dqoe_50;
input 	phy_ddio_dqoe_51;
input 	phy_ddio_dqs_dout_8;
input 	phy_ddio_dqs_dout_9;
input 	phy_ddio_dqs_dout_10;
input 	phy_ddio_dqs_dout_11;
input 	phy_ddio_dqslogic_aclr_fifoctrl_2;
input 	phy_ddio_dqslogic_aclr_pstamble_2;
input 	phy_ddio_dqslogic_dqsena_4;
input 	phy_ddio_dqslogic_dqsena_5;
input 	phy_ddio_dqslogic_fiforeset_2;
input 	phy_ddio_dqslogic_incrdataen_4;
input 	phy_ddio_dqslogic_incrdataen_5;
input 	phy_ddio_dqslogic_incwrptr_4;
input 	phy_ddio_dqslogic_incwrptr_5;
input 	phy_ddio_dqslogic_oct_4;
input 	phy_ddio_dqslogic_oct_5;
input 	phy_ddio_dqslogic_readlatency_10;
input 	phy_ddio_dqslogic_readlatency_11;
input 	phy_ddio_dqslogic_readlatency_12;
input 	phy_ddio_dqslogic_readlatency_13;
input 	phy_ddio_dqslogic_readlatency_14;
input 	phy_ddio_dqs_oe_4;
input 	phy_ddio_dqs_oe_5;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_11,phy_ddio_dmdout_10,phy_ddio_dmdout_9,phy_ddio_dmdout_8}),
	.write_data_in({phy_ddio_dqdout_103,phy_ddio_dqdout_102,phy_ddio_dqdout_101,phy_ddio_dqdout_100,phy_ddio_dqdout_99,phy_ddio_dqdout_98,phy_ddio_dqdout_97,phy_ddio_dqdout_96,phy_ddio_dqdout_95,phy_ddio_dqdout_94,phy_ddio_dqdout_93,phy_ddio_dqdout_92,phy_ddio_dqdout_91,phy_ddio_dqdout_90,
phy_ddio_dqdout_89,phy_ddio_dqdout_88,phy_ddio_dqdout_87,phy_ddio_dqdout_86,phy_ddio_dqdout_85,phy_ddio_dqdout_84,phy_ddio_dqdout_83,phy_ddio_dqdout_82,phy_ddio_dqdout_81,phy_ddio_dqdout_80,phy_ddio_dqdout_79,phy_ddio_dqdout_78,phy_ddio_dqdout_77,phy_ddio_dqdout_76,
phy_ddio_dqdout_75,phy_ddio_dqdout_74,phy_ddio_dqdout_73,phy_ddio_dqdout_72}),
	.write_oe_in({phy_ddio_dqoe_51,phy_ddio_dqoe_50,phy_ddio_dqoe_49,phy_ddio_dqoe_48,phy_ddio_dqoe_47,phy_ddio_dqoe_46,phy_ddio_dqoe_45,phy_ddio_dqoe_44,phy_ddio_dqoe_43,phy_ddio_dqoe_42,phy_ddio_dqoe_41,phy_ddio_dqoe_40,phy_ddio_dqoe_39,phy_ddio_dqoe_38,phy_ddio_dqoe_37,phy_ddio_dqoe_36}),
	.write_strobe({phy_ddio_dqs_dout_11,phy_ddio_dqs_dout_10,phy_ddio_dqs_dout_9,phy_ddio_dqs_dout_8}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_2),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_2),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_5,phy_ddio_dqslogic_dqsena_4}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_2),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_5,phy_ddio_dqslogic_incrdataen_4}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_5,phy_ddio_dqslogic_incwrptr_4}),
	.oct_ena_in({phy_ddio_dqslogic_oct_5,phy_ddio_dqslogic_oct_4}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_14,phy_ddio_dqslogic_readlatency_13,phy_ddio_dqslogic_readlatency_12,phy_ddio_dqslogic_readlatency_11,phy_ddio_dqslogic_readlatency_10}),
	.output_strobe_ena({phy_ddio_dqs_oe_5,phy_ddio_dqs_oe_4}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_2 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_altdqdqs_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	afi_clk,
	pll_write_clk,
	extra_output_pad_gen0delayed_data_out,
	phy_ddio_dmdout_12,
	phy_ddio_dmdout_13,
	phy_ddio_dmdout_14,
	phy_ddio_dmdout_15,
	phy_ddio_dqdout_108,
	phy_ddio_dqdout_109,
	phy_ddio_dqdout_110,
	phy_ddio_dqdout_111,
	phy_ddio_dqdout_112,
	phy_ddio_dqdout_113,
	phy_ddio_dqdout_114,
	phy_ddio_dqdout_115,
	phy_ddio_dqdout_116,
	phy_ddio_dqdout_117,
	phy_ddio_dqdout_118,
	phy_ddio_dqdout_119,
	phy_ddio_dqdout_120,
	phy_ddio_dqdout_121,
	phy_ddio_dqdout_122,
	phy_ddio_dqdout_123,
	phy_ddio_dqdout_124,
	phy_ddio_dqdout_125,
	phy_ddio_dqdout_126,
	phy_ddio_dqdout_127,
	phy_ddio_dqdout_128,
	phy_ddio_dqdout_129,
	phy_ddio_dqdout_130,
	phy_ddio_dqdout_131,
	phy_ddio_dqdout_132,
	phy_ddio_dqdout_133,
	phy_ddio_dqdout_134,
	phy_ddio_dqdout_135,
	phy_ddio_dqdout_136,
	phy_ddio_dqdout_137,
	phy_ddio_dqdout_138,
	phy_ddio_dqdout_139,
	phy_ddio_dqoe_54,
	phy_ddio_dqoe_55,
	phy_ddio_dqoe_56,
	phy_ddio_dqoe_57,
	phy_ddio_dqoe_58,
	phy_ddio_dqoe_59,
	phy_ddio_dqoe_60,
	phy_ddio_dqoe_61,
	phy_ddio_dqoe_62,
	phy_ddio_dqoe_63,
	phy_ddio_dqoe_64,
	phy_ddio_dqoe_65,
	phy_ddio_dqoe_66,
	phy_ddio_dqoe_67,
	phy_ddio_dqoe_68,
	phy_ddio_dqoe_69,
	phy_ddio_dqs_dout_12,
	phy_ddio_dqs_dout_13,
	phy_ddio_dqs_dout_14,
	phy_ddio_dqs_dout_15,
	phy_ddio_dqslogic_aclr_fifoctrl_3,
	phy_ddio_dqslogic_aclr_pstamble_3,
	phy_ddio_dqslogic_dqsena_6,
	phy_ddio_dqslogic_dqsena_7,
	phy_ddio_dqslogic_fiforeset_3,
	phy_ddio_dqslogic_incrdataen_6,
	phy_ddio_dqslogic_incrdataen_7,
	phy_ddio_dqslogic_incwrptr_6,
	phy_ddio_dqslogic_incwrptr_7,
	phy_ddio_dqslogic_oct_6,
	phy_ddio_dqslogic_oct_7,
	phy_ddio_dqslogic_readlatency_15,
	phy_ddio_dqslogic_readlatency_16,
	phy_ddio_dqslogic_readlatency_17,
	phy_ddio_dqslogic_readlatency_18,
	phy_ddio_dqslogic_readlatency_19,
	phy_ddio_dqs_oe_6,
	phy_ddio_dqs_oe_7,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	input_path_gen0read_fifo_out_0,
	input_path_gen0read_fifo_out_1,
	input_path_gen0read_fifo_out_2,
	input_path_gen0read_fifo_out_3,
	input_path_gen1read_fifo_out_0,
	input_path_gen1read_fifo_out_1,
	input_path_gen1read_fifo_out_2,
	input_path_gen1read_fifo_out_3,
	input_path_gen2read_fifo_out_0,
	input_path_gen2read_fifo_out_1,
	input_path_gen2read_fifo_out_2,
	input_path_gen2read_fifo_out_3,
	input_path_gen3read_fifo_out_0,
	input_path_gen3read_fifo_out_1,
	input_path_gen3read_fifo_out_2,
	input_path_gen3read_fifo_out_3,
	input_path_gen4read_fifo_out_0,
	input_path_gen4read_fifo_out_1,
	input_path_gen4read_fifo_out_2,
	input_path_gen4read_fifo_out_3,
	input_path_gen5read_fifo_out_0,
	input_path_gen5read_fifo_out_1,
	input_path_gen5read_fifo_out_2,
	input_path_gen5read_fifo_out_3,
	input_path_gen6read_fifo_out_0,
	input_path_gen6read_fifo_out_1,
	input_path_gen6read_fifo_out_2,
	input_path_gen6read_fifo_out_3,
	input_path_gen7read_fifo_out_0,
	input_path_gen7read_fifo_out_1,
	input_path_gen7read_fifo_out_2,
	input_path_gen7read_fifo_out_3,
	lfifo_rdata_valid,
	dll_delayctrl_0,
	dll_delayctrl_1,
	dll_delayctrl_2,
	dll_delayctrl_3,
	dll_delayctrl_4,
	dll_delayctrl_5,
	dll_delayctrl_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	afi_clk;
input 	pll_write_clk;
output 	extra_output_pad_gen0delayed_data_out;
input 	phy_ddio_dmdout_12;
input 	phy_ddio_dmdout_13;
input 	phy_ddio_dmdout_14;
input 	phy_ddio_dmdout_15;
input 	phy_ddio_dqdout_108;
input 	phy_ddio_dqdout_109;
input 	phy_ddio_dqdout_110;
input 	phy_ddio_dqdout_111;
input 	phy_ddio_dqdout_112;
input 	phy_ddio_dqdout_113;
input 	phy_ddio_dqdout_114;
input 	phy_ddio_dqdout_115;
input 	phy_ddio_dqdout_116;
input 	phy_ddio_dqdout_117;
input 	phy_ddio_dqdout_118;
input 	phy_ddio_dqdout_119;
input 	phy_ddio_dqdout_120;
input 	phy_ddio_dqdout_121;
input 	phy_ddio_dqdout_122;
input 	phy_ddio_dqdout_123;
input 	phy_ddio_dqdout_124;
input 	phy_ddio_dqdout_125;
input 	phy_ddio_dqdout_126;
input 	phy_ddio_dqdout_127;
input 	phy_ddio_dqdout_128;
input 	phy_ddio_dqdout_129;
input 	phy_ddio_dqdout_130;
input 	phy_ddio_dqdout_131;
input 	phy_ddio_dqdout_132;
input 	phy_ddio_dqdout_133;
input 	phy_ddio_dqdout_134;
input 	phy_ddio_dqdout_135;
input 	phy_ddio_dqdout_136;
input 	phy_ddio_dqdout_137;
input 	phy_ddio_dqdout_138;
input 	phy_ddio_dqdout_139;
input 	phy_ddio_dqoe_54;
input 	phy_ddio_dqoe_55;
input 	phy_ddio_dqoe_56;
input 	phy_ddio_dqoe_57;
input 	phy_ddio_dqoe_58;
input 	phy_ddio_dqoe_59;
input 	phy_ddio_dqoe_60;
input 	phy_ddio_dqoe_61;
input 	phy_ddio_dqoe_62;
input 	phy_ddio_dqoe_63;
input 	phy_ddio_dqoe_64;
input 	phy_ddio_dqoe_65;
input 	phy_ddio_dqoe_66;
input 	phy_ddio_dqoe_67;
input 	phy_ddio_dqoe_68;
input 	phy_ddio_dqoe_69;
input 	phy_ddio_dqs_dout_12;
input 	phy_ddio_dqs_dout_13;
input 	phy_ddio_dqs_dout_14;
input 	phy_ddio_dqs_dout_15;
input 	phy_ddio_dqslogic_aclr_fifoctrl_3;
input 	phy_ddio_dqslogic_aclr_pstamble_3;
input 	phy_ddio_dqslogic_dqsena_6;
input 	phy_ddio_dqslogic_dqsena_7;
input 	phy_ddio_dqslogic_fiforeset_3;
input 	phy_ddio_dqslogic_incrdataen_6;
input 	phy_ddio_dqslogic_incrdataen_7;
input 	phy_ddio_dqslogic_incwrptr_6;
input 	phy_ddio_dqslogic_incwrptr_7;
input 	phy_ddio_dqslogic_oct_6;
input 	phy_ddio_dqslogic_oct_7;
input 	phy_ddio_dqslogic_readlatency_15;
input 	phy_ddio_dqslogic_readlatency_16;
input 	phy_ddio_dqslogic_readlatency_17;
input 	phy_ddio_dqslogic_readlatency_18;
input 	phy_ddio_dqslogic_readlatency_19;
input 	phy_ddio_dqs_oe_6;
input 	phy_ddio_dqs_oe_7;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	input_path_gen0read_fifo_out_0;
output 	input_path_gen0read_fifo_out_1;
output 	input_path_gen0read_fifo_out_2;
output 	input_path_gen0read_fifo_out_3;
output 	input_path_gen1read_fifo_out_0;
output 	input_path_gen1read_fifo_out_1;
output 	input_path_gen1read_fifo_out_2;
output 	input_path_gen1read_fifo_out_3;
output 	input_path_gen2read_fifo_out_0;
output 	input_path_gen2read_fifo_out_1;
output 	input_path_gen2read_fifo_out_2;
output 	input_path_gen2read_fifo_out_3;
output 	input_path_gen3read_fifo_out_0;
output 	input_path_gen3read_fifo_out_1;
output 	input_path_gen3read_fifo_out_2;
output 	input_path_gen3read_fifo_out_3;
output 	input_path_gen4read_fifo_out_0;
output 	input_path_gen4read_fifo_out_1;
output 	input_path_gen4read_fifo_out_2;
output 	input_path_gen4read_fifo_out_3;
output 	input_path_gen5read_fifo_out_0;
output 	input_path_gen5read_fifo_out_1;
output 	input_path_gen5read_fifo_out_2;
output 	input_path_gen5read_fifo_out_3;
output 	input_path_gen6read_fifo_out_0;
output 	input_path_gen6read_fifo_out_1;
output 	input_path_gen6read_fifo_out_2;
output 	input_path_gen6read_fifo_out_3;
output 	input_path_gen7read_fifo_out_0;
output 	input_path_gen7read_fifo_out_1;
output 	input_path_gen7read_fifo_out_2;
output 	input_path_gen7read_fifo_out_3;
output 	lfifo_rdata_valid;
input 	dll_delayctrl_0;
input 	dll_delayctrl_1;
input 	dll_delayctrl_2;
input 	dll_delayctrl_3;
input 	dll_delayctrl_4;
input 	dll_delayctrl_5;
input 	dll_delayctrl_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 altdq_dqs2_inst(
	.dqsin(dqsin),
	.pad_gen0raw_input(pad_gen0raw_input),
	.pad_gen1raw_input(pad_gen1raw_input),
	.pad_gen2raw_input(pad_gen2raw_input),
	.pad_gen3raw_input(pad_gen3raw_input),
	.pad_gen4raw_input(pad_gen4raw_input),
	.pad_gen5raw_input(pad_gen5raw_input),
	.pad_gen6raw_input(pad_gen6raw_input),
	.pad_gen7raw_input(pad_gen7raw_input),
	.config_clock_in(afi_clk),
	.hr_clock_in(afi_clk),
	.write_strobe_clock_in(afi_clk),
	.fr_clock_in(pll_write_clk),
	.extra_output_pad_gen0delayed_data_out(extra_output_pad_gen0delayed_data_out),
	.extra_write_data_in({phy_ddio_dmdout_15,phy_ddio_dmdout_14,phy_ddio_dmdout_13,phy_ddio_dmdout_12}),
	.write_data_in({phy_ddio_dqdout_139,phy_ddio_dqdout_138,phy_ddio_dqdout_137,phy_ddio_dqdout_136,phy_ddio_dqdout_135,phy_ddio_dqdout_134,phy_ddio_dqdout_133,phy_ddio_dqdout_132,phy_ddio_dqdout_131,phy_ddio_dqdout_130,phy_ddio_dqdout_129,phy_ddio_dqdout_128,phy_ddio_dqdout_127,
phy_ddio_dqdout_126,phy_ddio_dqdout_125,phy_ddio_dqdout_124,phy_ddio_dqdout_123,phy_ddio_dqdout_122,phy_ddio_dqdout_121,phy_ddio_dqdout_120,phy_ddio_dqdout_119,phy_ddio_dqdout_118,phy_ddio_dqdout_117,phy_ddio_dqdout_116,phy_ddio_dqdout_115,phy_ddio_dqdout_114,
phy_ddio_dqdout_113,phy_ddio_dqdout_112,phy_ddio_dqdout_111,phy_ddio_dqdout_110,phy_ddio_dqdout_109,phy_ddio_dqdout_108}),
	.write_oe_in({phy_ddio_dqoe_69,phy_ddio_dqoe_68,phy_ddio_dqoe_67,phy_ddio_dqoe_66,phy_ddio_dqoe_65,phy_ddio_dqoe_64,phy_ddio_dqoe_63,phy_ddio_dqoe_62,phy_ddio_dqoe_61,phy_ddio_dqoe_60,phy_ddio_dqoe_59,phy_ddio_dqoe_58,phy_ddio_dqoe_57,phy_ddio_dqoe_56,phy_ddio_dqoe_55,phy_ddio_dqoe_54}),
	.write_strobe({phy_ddio_dqs_dout_15,phy_ddio_dqs_dout_14,phy_ddio_dqs_dout_13,phy_ddio_dqs_dout_12}),
	.lfifo_reset_n(phy_ddio_dqslogic_aclr_fifoctrl_3),
	.vfifo_reset_n(phy_ddio_dqslogic_aclr_pstamble_3),
	.lfifo_rdata_en_full({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.vfifo_qvld({phy_ddio_dqslogic_dqsena_7,phy_ddio_dqslogic_dqsena_6}),
	.rfifo_reset_n(phy_ddio_dqslogic_fiforeset_3),
	.lfifo_rdata_en({phy_ddio_dqslogic_incrdataen_7,phy_ddio_dqslogic_incrdataen_6}),
	.vfifo_inc_wr_ptr({phy_ddio_dqslogic_incwrptr_7,phy_ddio_dqslogic_incwrptr_6}),
	.oct_ena_in({phy_ddio_dqslogic_oct_7,phy_ddio_dqslogic_oct_6}),
	.lfifo_rd_latency({phy_ddio_dqslogic_readlatency_19,phy_ddio_dqslogic_readlatency_18,phy_ddio_dqslogic_readlatency_17,phy_ddio_dqslogic_readlatency_16,phy_ddio_dqslogic_readlatency_15}),
	.output_strobe_ena({phy_ddio_dqs_oe_7,phy_ddio_dqs_oe_6}),
	.pad_gen0delayed_data_out(pad_gen0delayed_data_out),
	.pad_gen0delayed_oe_1(pad_gen0delayed_oe_1),
	.delayed_oct(delayed_oct),
	.pad_gen1delayed_data_out(pad_gen1delayed_data_out),
	.pad_gen1delayed_oe_1(pad_gen1delayed_oe_1),
	.pad_gen2delayed_data_out(pad_gen2delayed_data_out),
	.pad_gen2delayed_oe_1(pad_gen2delayed_oe_1),
	.pad_gen3delayed_data_out(pad_gen3delayed_data_out),
	.pad_gen3delayed_oe_1(pad_gen3delayed_oe_1),
	.pad_gen4delayed_data_out(pad_gen4delayed_data_out),
	.pad_gen4delayed_oe_1(pad_gen4delayed_oe_1),
	.pad_gen5delayed_data_out(pad_gen5delayed_data_out),
	.pad_gen5delayed_oe_1(pad_gen5delayed_oe_1),
	.pad_gen6delayed_data_out(pad_gen6delayed_data_out),
	.pad_gen6delayed_oe_1(pad_gen6delayed_oe_1),
	.pad_gen7delayed_data_out(pad_gen7delayed_data_out),
	.pad_gen7delayed_oe_1(pad_gen7delayed_oe_1),
	.os(os),
	.os_bar(os_bar),
	.diff_oe(diff_oe),
	.diff_oe_bar(diff_oe_bar),
	.diff_dtc(diff_dtc),
	.diff_dtc_bar(diff_dtc_bar),
	.read_data_out({input_path_gen7read_fifo_out_3,input_path_gen7read_fifo_out_2,input_path_gen7read_fifo_out_1,input_path_gen7read_fifo_out_0,input_path_gen6read_fifo_out_3,input_path_gen6read_fifo_out_2,input_path_gen6read_fifo_out_1,input_path_gen6read_fifo_out_0,
input_path_gen5read_fifo_out_3,input_path_gen5read_fifo_out_2,input_path_gen5read_fifo_out_1,input_path_gen5read_fifo_out_0,input_path_gen4read_fifo_out_3,input_path_gen4read_fifo_out_2,input_path_gen4read_fifo_out_1,input_path_gen4read_fifo_out_0,
input_path_gen3read_fifo_out_3,input_path_gen3read_fifo_out_2,input_path_gen3read_fifo_out_1,input_path_gen3read_fifo_out_0,input_path_gen2read_fifo_out_3,input_path_gen2read_fifo_out_2,input_path_gen2read_fifo_out_1,input_path_gen2read_fifo_out_0,
input_path_gen1read_fifo_out_3,input_path_gen1read_fifo_out_2,input_path_gen1read_fifo_out_1,input_path_gen1read_fifo_out_0,input_path_gen0read_fifo_out_3,input_path_gen0read_fifo_out_2,input_path_gen0read_fifo_out_1,input_path_gen0read_fifo_out_0}),
	.lfifo_rdata_valid(lfifo_rdata_valid),
	.dll_delayctrl_in({dll_delayctrl_6,dll_delayctrl_5,dll_delayctrl_4,dll_delayctrl_3,dll_delayctrl_2,dll_delayctrl_1,dll_delayctrl_0}),
	.GND_port(GND_port));

endmodule

module terminal_qsys_altdq_dqs2_acv_connect_to_hard_phy_cyclonev_3 (
	dqsin,
	pad_gen0raw_input,
	pad_gen1raw_input,
	pad_gen2raw_input,
	pad_gen3raw_input,
	pad_gen4raw_input,
	pad_gen5raw_input,
	pad_gen6raw_input,
	pad_gen7raw_input,
	config_clock_in,
	hr_clock_in,
	write_strobe_clock_in,
	fr_clock_in,
	extra_output_pad_gen0delayed_data_out,
	extra_write_data_in,
	write_data_in,
	write_oe_in,
	write_strobe,
	lfifo_reset_n,
	vfifo_reset_n,
	lfifo_rdata_en_full,
	vfifo_qvld,
	rfifo_reset_n,
	lfifo_rdata_en,
	vfifo_inc_wr_ptr,
	oct_ena_in,
	lfifo_rd_latency,
	output_strobe_ena,
	pad_gen0delayed_data_out,
	pad_gen0delayed_oe_1,
	delayed_oct,
	pad_gen1delayed_data_out,
	pad_gen1delayed_oe_1,
	pad_gen2delayed_data_out,
	pad_gen2delayed_oe_1,
	pad_gen3delayed_data_out,
	pad_gen3delayed_oe_1,
	pad_gen4delayed_data_out,
	pad_gen4delayed_oe_1,
	pad_gen5delayed_data_out,
	pad_gen5delayed_oe_1,
	pad_gen6delayed_data_out,
	pad_gen6delayed_oe_1,
	pad_gen7delayed_data_out,
	pad_gen7delayed_oe_1,
	os,
	os_bar,
	diff_oe,
	diff_oe_bar,
	diff_dtc,
	diff_dtc_bar,
	read_data_out,
	lfifo_rdata_valid,
	dll_delayctrl_in,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	dqsin;
input 	pad_gen0raw_input;
input 	pad_gen1raw_input;
input 	pad_gen2raw_input;
input 	pad_gen3raw_input;
input 	pad_gen4raw_input;
input 	pad_gen5raw_input;
input 	pad_gen6raw_input;
input 	pad_gen7raw_input;
input 	config_clock_in;
input 	hr_clock_in;
input 	write_strobe_clock_in;
input 	fr_clock_in;
output 	extra_output_pad_gen0delayed_data_out;
input 	[3:0] extra_write_data_in;
input 	[31:0] write_data_in;
input 	[15:0] write_oe_in;
input 	[3:0] write_strobe;
input 	lfifo_reset_n;
input 	vfifo_reset_n;
input 	[1:0] lfifo_rdata_en_full;
input 	[1:0] vfifo_qvld;
input 	rfifo_reset_n;
input 	[1:0] lfifo_rdata_en;
input 	[1:0] vfifo_inc_wr_ptr;
input 	[1:0] oct_ena_in;
input 	[4:0] lfifo_rd_latency;
input 	[1:0] output_strobe_ena;
output 	pad_gen0delayed_data_out;
output 	pad_gen0delayed_oe_1;
output 	delayed_oct;
output 	pad_gen1delayed_data_out;
output 	pad_gen1delayed_oe_1;
output 	pad_gen2delayed_data_out;
output 	pad_gen2delayed_oe_1;
output 	pad_gen3delayed_data_out;
output 	pad_gen3delayed_oe_1;
output 	pad_gen4delayed_data_out;
output 	pad_gen4delayed_oe_1;
output 	pad_gen5delayed_data_out;
output 	pad_gen5delayed_oe_1;
output 	pad_gen6delayed_data_out;
output 	pad_gen6delayed_oe_1;
output 	pad_gen7delayed_data_out;
output 	pad_gen7delayed_oe_1;
output 	os;
output 	os_bar;
output 	diff_oe;
output 	diff_oe_bar;
output 	diff_dtc;
output 	diff_dtc_bar;
output 	[31:0] read_data_out;
output 	lfifo_rdata_valid;
input 	[6:0] dll_delayctrl_in;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \extra_output_pad_gen[0].config_1~dataout ;
wire \input_path_gen[0].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[1].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[2].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[3].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[4].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[5].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[6].read_fifo~O_LVDSMODEEN ;
wire \input_path_gen[7].read_fifo~O_LVDSMODEEN ;
wire \pad_gen[0].config_1~dataout ;
wire \dqs_config_gen[0].dqs_config_inst~dataout ;
wire \pad_gen[1].config_1~dataout ;
wire \pad_gen[2].config_1~dataout ;
wire \pad_gen[3].config_1~dataout ;
wire \pad_gen[4].config_1~dataout ;
wire \pad_gen[5].config_1~dataout ;
wire \pad_gen[6].config_1~dataout ;
wire \pad_gen[7].config_1~dataout ;
wire \leveled_dq_clocks[1] ;
wire \leveled_dq_clocks[2] ;
wire \leveled_dq_clocks[3] ;
wire \dqs_io_config_1~dataout ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;
wire lfifo_rden;
wire lfifo_oct;
wire \leveled_hr_clocks[0] ;
wire hr_seq_clock;
wire \extra_output_pad_gen[0].extra_outputhalfratebypass ;
wire \extra_output_pad_gen[0].fr_data_lo ;
wire \extra_output_pad_gen[0].fr_data_hi ;
wire \leveled_dq_clocks[0] ;
wire dq_shifted_clock;
wire \extra_output_pad_gen[0].aligned_data ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ;
wire \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ;
wire \dq_outputhalfratebypass[0] ;
wire \output_path_gen[0].fr_data_lo ;
wire \output_path_gen[0].fr_data_hi ;
wire \pad_gen[0].predelayed_data ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[0].fr_oe ;
wire \output_path_gen[0].oe_reg~q ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[0].dq_outputenabledelaysetting_dlc[4] ;
wire \dqshalfratebypass[0] ;
wire fr_os_oct;
wire \leveled_dqs_clocks[0] ;
wire dqs_shifted_clock;
wire predelayed_os_oct;
wire \octdelaysetting1_dlc[0][0] ;
wire \octdelaysetting1_dlc[0][1] ;
wire \octdelaysetting1_dlc[0][2] ;
wire \octdelaysetting1_dlc[0][3] ;
wire \octdelaysetting1_dlc[0][4] ;
wire \dq_outputhalfratebypass[1] ;
wire \output_path_gen[1].fr_data_lo ;
wire \output_path_gen[1].fr_data_hi ;
wire \pad_gen[1].predelayed_data ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[1].fr_oe ;
wire \output_path_gen[1].oe_reg~q ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[1].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[2] ;
wire \output_path_gen[2].fr_data_lo ;
wire \output_path_gen[2].fr_data_hi ;
wire \pad_gen[2].predelayed_data ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[2].fr_oe ;
wire \output_path_gen[2].oe_reg~q ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[2].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[3] ;
wire \output_path_gen[3].fr_data_lo ;
wire \output_path_gen[3].fr_data_hi ;
wire \pad_gen[3].predelayed_data ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[3].fr_oe ;
wire \output_path_gen[3].oe_reg~q ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[3].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[4] ;
wire \output_path_gen[4].fr_data_lo ;
wire \output_path_gen[4].fr_data_hi ;
wire \pad_gen[4].predelayed_data ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[4].fr_oe ;
wire \output_path_gen[4].oe_reg~q ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[4].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[5] ;
wire \output_path_gen[5].fr_data_lo ;
wire \output_path_gen[5].fr_data_hi ;
wire \pad_gen[5].predelayed_data ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[5].fr_oe ;
wire \output_path_gen[5].oe_reg~q ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[5].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[6] ;
wire \output_path_gen[6].fr_data_lo ;
wire \output_path_gen[6].fr_data_hi ;
wire \pad_gen[6].predelayed_data ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[6].fr_oe ;
wire \output_path_gen[6].oe_reg~q ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[6].dq_outputenabledelaysetting_dlc[4] ;
wire \dq_outputhalfratebypass[7] ;
wire \output_path_gen[7].fr_data_lo ;
wire \output_path_gen[7].fr_data_hi ;
wire \pad_gen[7].predelayed_data ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputdelaysetting_dlc[4] ;
wire \output_path_gen[7].fr_oe ;
wire \output_path_gen[7].oe_reg~q ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[0] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[1] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[2] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[3] ;
wire \pad_gen[7].dq_outputenabledelaysetting_dlc[4] ;
wire fr_os_lo;
wire fr_os_hi;
wire predelayed_os;
wire \dqs_outputdelaysetting_dlc[0] ;
wire \dqs_outputdelaysetting_dlc[1] ;
wire \dqs_outputdelaysetting_dlc[2] ;
wire \dqs_outputdelaysetting_dlc[3] ;
wire \dqs_outputdelaysetting_dlc[4] ;
wire os_delayed2;
wire fr_os_oe;
wire \os_oe_reg~q ;
wire \dqs_outputenabledelaysetting_dlc[0] ;
wire \dqs_outputenabledelaysetting_dlc[1] ;
wire \dqs_outputenabledelaysetting_dlc[2] ;
wire \dqs_outputenabledelaysetting_dlc[3] ;
wire \dqs_outputenabledelaysetting_dlc[4] ;
wire delayed_os_oe;
wire \rfifo_clock_select[0] ;
wire \rfifo_clock_select[1] ;
wire \input_path_gen[0].rfifo_rd_clk ;
wire vfifo_inc_wr_ptr_fr;
wire vfifo_qvld_fr;
wire ena_zero_phase_clock;
wire dqs_pre_delayed;
wire \enadqsenablephasetransferreg[0] ;
wire \dqsenablectrlphaseinvert[0] ;
wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \dqsenablectrlphasesetting[0][0] ;
wire \dqsenablectrlphasesetting[0][1] ;
wire ena_clock;
wire dqs_enable_shifted;
wire \dqsenabledelaysetting_dlc[0][0] ;
wire \dqsenabledelaysetting_dlc[0][1] ;
wire \dqsenabledelaysetting_dlc[0][2] ;
wire \dqsenabledelaysetting_dlc[0][3] ;
wire \dqsenabledelaysetting_dlc[0][4] ;
wire dqs_enable_int;
wire \dqsdisabledelaysetting_dlc[0][0] ;
wire \dqsdisabledelaysetting_dlc[0][1] ;
wire \dqsdisabledelaysetting_dlc[0][2] ;
wire \dqsdisabledelaysetting_dlc[0][3] ;
wire \dqsdisabledelaysetting_dlc[0][4] ;
wire dqs_disable_int;
wire dqs_shifted;
wire \dqsbusoutdelaysetting_dlc[0][0] ;
wire \dqsbusoutdelaysetting_dlc[0][1] ;
wire \dqsbusoutdelaysetting_dlc[0][2] ;
wire \dqsbusoutdelaysetting_dlc[0][3] ;
wire \dqsbusoutdelaysetting_dlc[0][4] ;
wire dqsbusout;
wire \pad_gen[0].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[0].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[0] ;
wire \input_path_gen[0].aligned_input[0] ;
wire \input_path_gen[0].aligned_input[1] ;
wire \rfifo_mode[0] ;
wire \rfifo_mode[1] ;
wire \rfifo_mode[2] ;
wire \rfifo_clock_select[2] ;
wire \rfifo_clock_select[3] ;
wire \input_path_gen[1].rfifo_rd_clk ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[1].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[1] ;
wire \input_path_gen[1].aligned_input[0] ;
wire \input_path_gen[1].aligned_input[1] ;
wire \rfifo_mode[3] ;
wire \rfifo_mode[4] ;
wire \rfifo_mode[5] ;
wire \rfifo_clock_select[4] ;
wire \rfifo_clock_select[5] ;
wire \input_path_gen[2].rfifo_rd_clk ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[2].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[2] ;
wire \input_path_gen[2].aligned_input[0] ;
wire \input_path_gen[2].aligned_input[1] ;
wire \rfifo_mode[6] ;
wire \rfifo_mode[7] ;
wire \rfifo_mode[8] ;
wire \rfifo_clock_select[6] ;
wire \rfifo_clock_select[7] ;
wire \input_path_gen[3].rfifo_rd_clk ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[3].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[3] ;
wire \input_path_gen[3].aligned_input[0] ;
wire \input_path_gen[3].aligned_input[1] ;
wire \rfifo_mode[9] ;
wire \rfifo_mode[10] ;
wire \rfifo_mode[11] ;
wire \rfifo_clock_select[8] ;
wire \rfifo_clock_select[9] ;
wire \input_path_gen[4].rfifo_rd_clk ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[4].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[4] ;
wire \input_path_gen[4].aligned_input[0] ;
wire \input_path_gen[4].aligned_input[1] ;
wire \rfifo_mode[12] ;
wire \rfifo_mode[13] ;
wire \rfifo_mode[14] ;
wire \rfifo_clock_select[10] ;
wire \rfifo_clock_select[11] ;
wire \input_path_gen[5].rfifo_rd_clk ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[5].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[5] ;
wire \input_path_gen[5].aligned_input[0] ;
wire \input_path_gen[5].aligned_input[1] ;
wire \rfifo_mode[15] ;
wire \rfifo_mode[16] ;
wire \rfifo_mode[17] ;
wire \rfifo_clock_select[12] ;
wire \rfifo_clock_select[13] ;
wire \input_path_gen[6].rfifo_rd_clk ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[6].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[6] ;
wire \input_path_gen[6].aligned_input[0] ;
wire \input_path_gen[6].aligned_input[1] ;
wire \rfifo_mode[18] ;
wire \rfifo_mode[19] ;
wire \rfifo_mode[20] ;
wire \rfifo_clock_select[14] ;
wire \rfifo_clock_select[15] ;
wire \input_path_gen[7].rfifo_rd_clk ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[0] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[1] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[2] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[3] ;
wire \pad_gen[7].dq_inputdelaysetting_dlc[4] ;
wire \ddr_data[7] ;
wire \input_path_gen[7].aligned_input[0] ;
wire \input_path_gen[7].aligned_input[1] ;
wire \rfifo_mode[21] ;
wire \rfifo_mode[22] ;
wire \rfifo_mode[23] ;
wire lfifo_rdata_en_fr;
wire lfifo_rdata_en_full_fr;

wire [4:0] \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [3:0] \input_path_gen[0].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[1].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[2].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[3].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[4].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[5].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[6].read_fifo_DOUT_bus ;
wire [3:0] \input_path_gen[7].read_fifo_DOUT_bus ;
wire [4:0] \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[0].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ;
wire [1:0] \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ;
wire [4:0] \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[1].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[2].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[3].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[4].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[5].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[6].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [4:0] \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ;
wire [2:0] \pad_gen[7].config_1_READFIFOMODE_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ;
wire [4:0] \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ;
wire [1:0] \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ;
wire [3:0] leveling_delay_chain_dq_CLKOUT_bus;
wire [4:0] dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus;
wire [4:0] dqs_io_config_1_OUTPUTREGDELAYSETTING_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;
wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;

assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4]  = \extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign read_data_out[0] = \input_path_gen[0].read_fifo_DOUT_bus [0];
assign read_data_out[1] = \input_path_gen[0].read_fifo_DOUT_bus [1];
assign read_data_out[2] = \input_path_gen[0].read_fifo_DOUT_bus [2];
assign read_data_out[3] = \input_path_gen[0].read_fifo_DOUT_bus [3];

assign read_data_out[4] = \input_path_gen[1].read_fifo_DOUT_bus [0];
assign read_data_out[5] = \input_path_gen[1].read_fifo_DOUT_bus [1];
assign read_data_out[6] = \input_path_gen[1].read_fifo_DOUT_bus [2];
assign read_data_out[7] = \input_path_gen[1].read_fifo_DOUT_bus [3];

assign read_data_out[8] = \input_path_gen[2].read_fifo_DOUT_bus [0];
assign read_data_out[9] = \input_path_gen[2].read_fifo_DOUT_bus [1];
assign read_data_out[10] = \input_path_gen[2].read_fifo_DOUT_bus [2];
assign read_data_out[11] = \input_path_gen[2].read_fifo_DOUT_bus [3];

assign read_data_out[12] = \input_path_gen[3].read_fifo_DOUT_bus [0];
assign read_data_out[13] = \input_path_gen[3].read_fifo_DOUT_bus [1];
assign read_data_out[14] = \input_path_gen[3].read_fifo_DOUT_bus [2];
assign read_data_out[15] = \input_path_gen[3].read_fifo_DOUT_bus [3];

assign read_data_out[16] = \input_path_gen[4].read_fifo_DOUT_bus [0];
assign read_data_out[17] = \input_path_gen[4].read_fifo_DOUT_bus [1];
assign read_data_out[18] = \input_path_gen[4].read_fifo_DOUT_bus [2];
assign read_data_out[19] = \input_path_gen[4].read_fifo_DOUT_bus [3];

assign read_data_out[20] = \input_path_gen[5].read_fifo_DOUT_bus [0];
assign read_data_out[21] = \input_path_gen[5].read_fifo_DOUT_bus [1];
assign read_data_out[22] = \input_path_gen[5].read_fifo_DOUT_bus [2];
assign read_data_out[23] = \input_path_gen[5].read_fifo_DOUT_bus [3];

assign read_data_out[24] = \input_path_gen[6].read_fifo_DOUT_bus [0];
assign read_data_out[25] = \input_path_gen[6].read_fifo_DOUT_bus [1];
assign read_data_out[26] = \input_path_gen[6].read_fifo_DOUT_bus [2];
assign read_data_out[27] = \input_path_gen[6].read_fifo_DOUT_bus [3];

assign read_data_out[28] = \input_path_gen[7].read_fifo_DOUT_bus [0];
assign read_data_out[29] = \input_path_gen[7].read_fifo_DOUT_bus [1];
assign read_data_out[30] = \input_path_gen[7].read_fifo_DOUT_bus [2];
assign read_data_out[31] = \input_path_gen[7].read_fifo_DOUT_bus [3];

assign \pad_gen[0].dq_inputdelaysetting_dlc[0]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[0].dq_inputdelaysetting_dlc[1]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[0].dq_inputdelaysetting_dlc[2]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[0].dq_inputdelaysetting_dlc[3]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[0].dq_inputdelaysetting_dlc[4]  = \pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[0]  = \pad_gen[0].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[1]  = \pad_gen[0].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[2]  = \pad_gen[0].config_1_READFIFOMODE_bus [2];

assign \pad_gen[0].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[0].dq_outputdelaysetting_dlc[0]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[0].dq_outputdelaysetting_dlc[1]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[0].dq_outputdelaysetting_dlc[2]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[0].dq_outputdelaysetting_dlc[3]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[0].dq_outputdelaysetting_dlc[4]  = \pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[0]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[1]  = \pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \dqsbusoutdelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [0];
assign \dqsbusoutdelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [1];
assign \dqsbusoutdelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [2];
assign \dqsbusoutdelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [3];
assign \dqsbusoutdelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus [4];

assign \dqsenablectrlphasesetting[0][0]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [0];
assign \dqsenablectrlphasesetting[0][1]  = \dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus [1];

assign \octdelaysetting1_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [0];
assign \octdelaysetting1_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [1];
assign \octdelaysetting1_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [2];
assign \octdelaysetting1_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [3];
assign \octdelaysetting1_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus [4];

assign \dqsenabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [0];
assign \dqsenabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [1];
assign \dqsenabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [2];
assign \dqsenabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [3];
assign \dqsenabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus [4];

assign \dqsdisabledelaysetting_dlc[0][0]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [0];
assign \dqsdisabledelaysetting_dlc[0][1]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [1];
assign \dqsdisabledelaysetting_dlc[0][2]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [2];
assign \dqsdisabledelaysetting_dlc[0][3]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [3];
assign \dqsdisabledelaysetting_dlc[0][4]  = \dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus [4];

assign \pad_gen[1].dq_inputdelaysetting_dlc[0]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[1].dq_inputdelaysetting_dlc[1]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[1].dq_inputdelaysetting_dlc[2]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[1].dq_inputdelaysetting_dlc[3]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[1].dq_inputdelaysetting_dlc[4]  = \pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[3]  = \pad_gen[1].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[4]  = \pad_gen[1].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[5]  = \pad_gen[1].config_1_READFIFOMODE_bus [2];

assign \pad_gen[1].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[1].dq_outputdelaysetting_dlc[0]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[1].dq_outputdelaysetting_dlc[1]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[1].dq_outputdelaysetting_dlc[2]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[1].dq_outputdelaysetting_dlc[3]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[1].dq_outputdelaysetting_dlc[4]  = \pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[2]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[3]  = \pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[2].dq_inputdelaysetting_dlc[0]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[2].dq_inputdelaysetting_dlc[1]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[2].dq_inputdelaysetting_dlc[2]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[2].dq_inputdelaysetting_dlc[3]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[2].dq_inputdelaysetting_dlc[4]  = \pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[6]  = \pad_gen[2].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[7]  = \pad_gen[2].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[8]  = \pad_gen[2].config_1_READFIFOMODE_bus [2];

assign \pad_gen[2].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[2].dq_outputdelaysetting_dlc[0]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[2].dq_outputdelaysetting_dlc[1]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[2].dq_outputdelaysetting_dlc[2]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[2].dq_outputdelaysetting_dlc[3]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[2].dq_outputdelaysetting_dlc[4]  = \pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[4]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[5]  = \pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[3].dq_inputdelaysetting_dlc[0]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[3].dq_inputdelaysetting_dlc[1]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[3].dq_inputdelaysetting_dlc[2]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[3].dq_inputdelaysetting_dlc[3]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[3].dq_inputdelaysetting_dlc[4]  = \pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[9]  = \pad_gen[3].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[10]  = \pad_gen[3].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[11]  = \pad_gen[3].config_1_READFIFOMODE_bus [2];

assign \pad_gen[3].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[3].dq_outputdelaysetting_dlc[0]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[3].dq_outputdelaysetting_dlc[1]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[3].dq_outputdelaysetting_dlc[2]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[3].dq_outputdelaysetting_dlc[3]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[3].dq_outputdelaysetting_dlc[4]  = \pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[6]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[7]  = \pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[4].dq_inputdelaysetting_dlc[0]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[4].dq_inputdelaysetting_dlc[1]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[4].dq_inputdelaysetting_dlc[2]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[4].dq_inputdelaysetting_dlc[3]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[4].dq_inputdelaysetting_dlc[4]  = \pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[12]  = \pad_gen[4].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[13]  = \pad_gen[4].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[14]  = \pad_gen[4].config_1_READFIFOMODE_bus [2];

assign \pad_gen[4].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[4].dq_outputdelaysetting_dlc[0]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[4].dq_outputdelaysetting_dlc[1]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[4].dq_outputdelaysetting_dlc[2]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[4].dq_outputdelaysetting_dlc[3]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[4].dq_outputdelaysetting_dlc[4]  = \pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[8]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[9]  = \pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[5].dq_inputdelaysetting_dlc[0]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[5].dq_inputdelaysetting_dlc[1]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[5].dq_inputdelaysetting_dlc[2]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[5].dq_inputdelaysetting_dlc[3]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[5].dq_inputdelaysetting_dlc[4]  = \pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[15]  = \pad_gen[5].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[16]  = \pad_gen[5].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[17]  = \pad_gen[5].config_1_READFIFOMODE_bus [2];

assign \pad_gen[5].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[5].dq_outputdelaysetting_dlc[0]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[5].dq_outputdelaysetting_dlc[1]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[5].dq_outputdelaysetting_dlc[2]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[5].dq_outputdelaysetting_dlc[3]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[5].dq_outputdelaysetting_dlc[4]  = \pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[10]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[11]  = \pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[6].dq_inputdelaysetting_dlc[0]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[6].dq_inputdelaysetting_dlc[1]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[6].dq_inputdelaysetting_dlc[2]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[6].dq_inputdelaysetting_dlc[3]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[6].dq_inputdelaysetting_dlc[4]  = \pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[18]  = \pad_gen[6].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[19]  = \pad_gen[6].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[20]  = \pad_gen[6].config_1_READFIFOMODE_bus [2];

assign \pad_gen[6].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[6].dq_outputdelaysetting_dlc[0]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[6].dq_outputdelaysetting_dlc[1]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[6].dq_outputdelaysetting_dlc[2]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[6].dq_outputdelaysetting_dlc[3]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[6].dq_outputdelaysetting_dlc[4]  = \pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[12]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[13]  = \pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \pad_gen[7].dq_inputdelaysetting_dlc[0]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [0];
assign \pad_gen[7].dq_inputdelaysetting_dlc[1]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [1];
assign \pad_gen[7].dq_inputdelaysetting_dlc[2]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [2];
assign \pad_gen[7].dq_inputdelaysetting_dlc[3]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [3];
assign \pad_gen[7].dq_inputdelaysetting_dlc[4]  = \pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus [4];

assign \rfifo_mode[21]  = \pad_gen[7].config_1_READFIFOMODE_bus [0];
assign \rfifo_mode[22]  = \pad_gen[7].config_1_READFIFOMODE_bus [1];
assign \rfifo_mode[23]  = \pad_gen[7].config_1_READFIFOMODE_bus [2];

assign \pad_gen[7].dq_outputenabledelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputenabledelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus [4];

assign \pad_gen[7].dq_outputdelaysetting_dlc[0]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [0];
assign \pad_gen[7].dq_outputdelaysetting_dlc[1]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [1];
assign \pad_gen[7].dq_outputdelaysetting_dlc[2]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [2];
assign \pad_gen[7].dq_outputdelaysetting_dlc[3]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [3];
assign \pad_gen[7].dq_outputdelaysetting_dlc[4]  = \pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus [4];

assign \rfifo_clock_select[14]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [0];
assign \rfifo_clock_select[15]  = \pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus [1];

assign \leveled_dq_clocks[0]  = leveling_delay_chain_dq_CLKOUT_bus[0];
assign \leveled_dq_clocks[1]  = leveling_delay_chain_dq_CLKOUT_bus[1];
assign \leveled_dq_clocks[2]  = leveling_delay_chain_dq_CLKOUT_bus[2];
assign \leveled_dq_clocks[3]  = leveling_delay_chain_dq_CLKOUT_bus[3];

assign \dqs_outputenabledelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[0];
assign \dqs_outputenabledelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[1];
assign \dqs_outputenabledelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[2];
assign \dqs_outputenabledelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[3];
assign \dqs_outputenabledelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus[4];

assign \dqs_outputdelaysetting_dlc[0]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[0];
assign \dqs_outputdelaysetting_dlc[1]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[1];
assign \dqs_outputdelaysetting_dlc[2]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[2];
assign \dqs_outputdelaysetting_dlc[3]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[3];
assign \dqs_outputdelaysetting_dlc[4]  = dqs_io_config_1_OUTPUTREGDELAYSETTING_bus[4];

assign \leveled_hr_clocks[0]  = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

assign \leveled_dqs_clocks[0]  = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

cyclonev_delay_chain \extra_output_pad_gen[0].out_delay_1 (
	.datain(\extra_output_pad_gen[0].aligned_data ),
	.delayctrlin({\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[4] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[3] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[2] ,\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[1] ,
\extra_output_pad_gen[0].dq_outputdelaysetting1_dlc[0] }),
	.dataout(extra_output_pad_gen0delayed_data_out));
defparam \extra_output_pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \extra_output_pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].out_delay_1 (
	.datain(\pad_gen[0].predelayed_data ),
	.delayctrlin({\pad_gen[0].dq_outputdelaysetting_dlc[4] ,\pad_gen[0].dq_outputdelaysetting_dlc[3] ,\pad_gen[0].dq_outputdelaysetting_dlc[2] ,\pad_gen[0].dq_outputdelaysetting_dlc[1] ,\pad_gen[0].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_data_out));
defparam \pad_gen[0].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].oe_delay_1 (
	.datain(\output_path_gen[0].oe_reg~q ),
	.delayctrlin({\pad_gen[0].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[0].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen0delayed_oe_1));
defparam \pad_gen[0].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[0].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain oct_delay(
	.datain(predelayed_os_oct),
	.delayctrlin({\octdelaysetting1_dlc[0][4] ,\octdelaysetting1_dlc[0][3] ,\octdelaysetting1_dlc[0][2] ,\octdelaysetting1_dlc[0][1] ,\octdelaysetting1_dlc[0][0] }),
	.dataout(delayed_oct));
defparam oct_delay.sim_falling_delay_increment = 10;
defparam oct_delay.sim_intrinsic_falling_delay = 0;
defparam oct_delay.sim_intrinsic_rising_delay = 0;
defparam oct_delay.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].out_delay_1 (
	.datain(\pad_gen[1].predelayed_data ),
	.delayctrlin({\pad_gen[1].dq_outputdelaysetting_dlc[4] ,\pad_gen[1].dq_outputdelaysetting_dlc[3] ,\pad_gen[1].dq_outputdelaysetting_dlc[2] ,\pad_gen[1].dq_outputdelaysetting_dlc[1] ,\pad_gen[1].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_data_out));
defparam \pad_gen[1].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[1].oe_delay_1 (
	.datain(\output_path_gen[1].oe_reg~q ),
	.delayctrlin({\pad_gen[1].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[1].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen1delayed_oe_1));
defparam \pad_gen[1].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[1].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].out_delay_1 (
	.datain(\pad_gen[2].predelayed_data ),
	.delayctrlin({\pad_gen[2].dq_outputdelaysetting_dlc[4] ,\pad_gen[2].dq_outputdelaysetting_dlc[3] ,\pad_gen[2].dq_outputdelaysetting_dlc[2] ,\pad_gen[2].dq_outputdelaysetting_dlc[1] ,\pad_gen[2].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_data_out));
defparam \pad_gen[2].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[2].oe_delay_1 (
	.datain(\output_path_gen[2].oe_reg~q ),
	.delayctrlin({\pad_gen[2].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[2].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen2delayed_oe_1));
defparam \pad_gen[2].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[2].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].out_delay_1 (
	.datain(\pad_gen[3].predelayed_data ),
	.delayctrlin({\pad_gen[3].dq_outputdelaysetting_dlc[4] ,\pad_gen[3].dq_outputdelaysetting_dlc[3] ,\pad_gen[3].dq_outputdelaysetting_dlc[2] ,\pad_gen[3].dq_outputdelaysetting_dlc[1] ,\pad_gen[3].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_data_out));
defparam \pad_gen[3].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[3].oe_delay_1 (
	.datain(\output_path_gen[3].oe_reg~q ),
	.delayctrlin({\pad_gen[3].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[3].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen3delayed_oe_1));
defparam \pad_gen[3].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[3].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].out_delay_1 (
	.datain(\pad_gen[4].predelayed_data ),
	.delayctrlin({\pad_gen[4].dq_outputdelaysetting_dlc[4] ,\pad_gen[4].dq_outputdelaysetting_dlc[3] ,\pad_gen[4].dq_outputdelaysetting_dlc[2] ,\pad_gen[4].dq_outputdelaysetting_dlc[1] ,\pad_gen[4].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_data_out));
defparam \pad_gen[4].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[4].oe_delay_1 (
	.datain(\output_path_gen[4].oe_reg~q ),
	.delayctrlin({\pad_gen[4].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[4].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen4delayed_oe_1));
defparam \pad_gen[4].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[4].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].out_delay_1 (
	.datain(\pad_gen[5].predelayed_data ),
	.delayctrlin({\pad_gen[5].dq_outputdelaysetting_dlc[4] ,\pad_gen[5].dq_outputdelaysetting_dlc[3] ,\pad_gen[5].dq_outputdelaysetting_dlc[2] ,\pad_gen[5].dq_outputdelaysetting_dlc[1] ,\pad_gen[5].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_data_out));
defparam \pad_gen[5].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[5].oe_delay_1 (
	.datain(\output_path_gen[5].oe_reg~q ),
	.delayctrlin({\pad_gen[5].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[5].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen5delayed_oe_1));
defparam \pad_gen[5].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[5].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].out_delay_1 (
	.datain(\pad_gen[6].predelayed_data ),
	.delayctrlin({\pad_gen[6].dq_outputdelaysetting_dlc[4] ,\pad_gen[6].dq_outputdelaysetting_dlc[3] ,\pad_gen[6].dq_outputdelaysetting_dlc[2] ,\pad_gen[6].dq_outputdelaysetting_dlc[1] ,\pad_gen[6].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_data_out));
defparam \pad_gen[6].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[6].oe_delay_1 (
	.datain(\output_path_gen[6].oe_reg~q ),
	.delayctrlin({\pad_gen[6].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[6].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen6delayed_oe_1));
defparam \pad_gen[6].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[6].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].out_delay_1 (
	.datain(\pad_gen[7].predelayed_data ),
	.delayctrlin({\pad_gen[7].dq_outputdelaysetting_dlc[4] ,\pad_gen[7].dq_outputdelaysetting_dlc[3] ,\pad_gen[7].dq_outputdelaysetting_dlc[2] ,\pad_gen[7].dq_outputdelaysetting_dlc[1] ,\pad_gen[7].dq_outputdelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_data_out));
defparam \pad_gen[7].out_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].out_delay_1 .sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[7].oe_delay_1 (
	.datain(\output_path_gen[7].oe_reg~q ),
	.delayctrlin({\pad_gen[7].dq_outputenabledelaysetting_dlc[4] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[3] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[2] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[1] ,\pad_gen[7].dq_outputenabledelaysetting_dlc[0] }),
	.dataout(pad_gen7delayed_oe_1));
defparam \pad_gen[7].oe_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_falling_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_intrinsic_rising_delay = 0;
defparam \pad_gen[7].oe_delay_1 .sim_rising_delay_increment = 10;

cyclonev_pseudo_diff_out pseudo_diffa_0(
	.i(os_delayed2),
	.oein(delayed_os_oe),
	.dtcin(delayed_oct),
	.o(os),
	.obar(os_bar),
	.oeout(diff_oe),
	.oebout(diff_oe_bar),
	.dtc(diff_dtc),
	.dtcbar(diff_dtc_bar));

cyclonev_ir_fifo_userdes \input_path_gen[0].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[0].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[0].aligned_input[1] ,\input_path_gen[0].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[2] ,\rfifo_mode[1] ,\rfifo_mode[0] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[0].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[0].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[0].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[0].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[0].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[0].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[0].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[0].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[0].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[0].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[1].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[1].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[1].aligned_input[1] ,\input_path_gen[1].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[5] ,\rfifo_mode[4] ,\rfifo_mode[3] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[1].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[1].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[1].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[1].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[1].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[1].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[1].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[1].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[1].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[1].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[2].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[2].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[2].aligned_input[1] ,\input_path_gen[2].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[8] ,\rfifo_mode[7] ,\rfifo_mode[6] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[2].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[2].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[2].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[2].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[2].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[2].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[2].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[2].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[2].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[2].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[3].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[3].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[3].aligned_input[1] ,\input_path_gen[3].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[11] ,\rfifo_mode[10] ,\rfifo_mode[9] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[3].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[3].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[3].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[3].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[3].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[3].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[3].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[3].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[3].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[3].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[4].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[4].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[4].aligned_input[1] ,\input_path_gen[4].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[14] ,\rfifo_mode[13] ,\rfifo_mode[12] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[4].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[4].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[4].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[4].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[4].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[4].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[4].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[4].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[4].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[4].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[5].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[5].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[5].aligned_input[1] ,\input_path_gen[5].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[17] ,\rfifo_mode[16] ,\rfifo_mode[15] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[5].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[5].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[5].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[5].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[5].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[5].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[5].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[5].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[5].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[5].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[6].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[6].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[6].aligned_input[1] ,\input_path_gen[6].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[20] ,\rfifo_mode[19] ,\rfifo_mode[18] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[6].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[6].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[6].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[6].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[6].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[6].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[6].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[6].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[6].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[6].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_ir_fifo_userdes \input_path_gen[7].read_fifo (
	.bslipctl(gnd),
	.bslipin(gnd),
	.loaden(gnd),
	.readclk(\input_path_gen[7].rfifo_rd_clk ),
	.readenable(lfifo_rden),
	.regscan(gnd),
	.regscanovrd(gnd),
	.rstn(rfifo_reset_n),
	.scanin(gnd),
	.tstclk(gnd),
	.writeclk(!dqsbusout),
	.writeenable(vcc),
	.dinfiforx({\input_path_gen[7].aligned_input[1] ,\input_path_gen[7].aligned_input[0] }),
	.dynfifomode({\rfifo_mode[23] ,\rfifo_mode[22] ,\rfifo_mode[21] }),
	.txin(10'b0000000000),
	.bslipmax(),
	.bslipout(),
	.lvdsmodeen(\input_path_gen[7].read_fifo~O_LVDSMODEEN ),
	.lvdstxsel(),
	.scanout(),
	.txout(),
	.dout(\input_path_gen[7].read_fifo_DOUT_bus ),
	.rxout());
defparam \input_path_gen[7].read_fifo .a_enable_soft_cdr = "false";
defparam \input_path_gen[7].read_fifo .a_rb_bslipcfg = 1;
defparam \input_path_gen[7].read_fifo .a_rb_bypass_serializer = "false";
defparam \input_path_gen[7].read_fifo .a_rb_data_width = 10;
defparam \input_path_gen[7].read_fifo .a_rb_fifo_mode = "hrate_mode";
defparam \input_path_gen[7].read_fifo .a_rb_tx_outclk = "false";
defparam \input_path_gen[7].read_fifo .a_sim_readenable_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_sim_wclk_pre_delay = 10;
defparam \input_path_gen[7].read_fifo .a_use_dynamic_fifo_mode = "true";

cyclonev_lfifo lfifo(
	.rdataen(lfifo_rdata_en_fr),
	.rdataenfull(lfifo_rdata_en_full_fr),
	.rstn(lfifo_reset_n),
	.clk(dqs_shifted_clock),
	.rdlatency({lfifo_rd_latency[4],lfifo_rd_latency[3],lfifo_rd_latency[2],lfifo_rd_latency[1],lfifo_rd_latency[0]}),
	.rdatavalid(lfifo_rdata_valid),
	.rden(lfifo_rden),
	.octlfifo(lfifo_oct));
defparam lfifo.oct_lfifo_enable = -1;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(config_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_hr(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_hr_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(hr_seq_clock));
defparam clk_phase_select_hr.invert_phase = "false";
defparam clk_phase_select_hr.phase_setting = 0;
defparam clk_phase_select_hr.physical_clock_source = "hr";
defparam clk_phase_select_hr.use_dqs_input = "false";
defparam clk_phase_select_hr.use_phasectrlin = "false";

cyclonev_io_config \extra_output_pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.dataout(\extra_output_pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(\extra_output_pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(),
	.padtoinputregisterdelaysetting());

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_lo (
	.datainlo(extra_write_data_in[3]),
	.datainhi(extra_write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \extra_output_pad_gen[0].hr_to_fr_hi (
	.datainlo(extra_write_data_in[2]),
	.datainhi(extra_write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\extra_output_pad_gen[0].extra_outputhalfratebypass ),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .power_up = "low";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \extra_output_pad_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dq(
	.clkin(fr_clock_in),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_dq_CLKOUT_bus));
defparam leveling_delay_chain_dq.physical_clock_source = "dq";
defparam leveling_delay_chain_dq.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dq.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dq(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dq_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dq_shifted_clock));
defparam clk_phase_select_dq.invert_phase = "false";
defparam clk_phase_select_dq.phase_setting = 0;
defparam clk_phase_select_dq.physical_clock_source = "dq";
defparam clk_phase_select_dq.use_dqs_input = "false";
defparam clk_phase_select_dq.use_phasectrlin = "false";

cyclonev_ddio_out \extra_output_pad_gen[0].ddio_out (
	.datainlo(\extra_output_pad_gen[0].fr_data_lo ),
	.datainhi(\extra_output_pad_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\extra_output_pad_gen[0].aligned_data ),
	.dfflo(),
	.dffhi());
defparam \extra_output_pad_gen[0].ddio_out .async_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .half_rate_mode = "false";
defparam \extra_output_pad_gen[0].ddio_out .power_up = "low";
defparam \extra_output_pad_gen[0].ddio_out .sync_mode = "none";
defparam \extra_output_pad_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_io_config \pad_gen[0].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[0] ),
	.dataout(\pad_gen[0].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[0].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[0].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[0].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[0].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[0].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_lo (
	.datainlo(write_data_in[3]),
	.datainhi(write_data_in[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_hi (
	.datainlo(write_data_in[2]),
	.datainhi(write_data_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].ddio_out (
	.datainlo(\output_path_gen[0].fr_data_lo ),
	.datainhi(\output_path_gen[0].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[0].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].ddio_out .async_mode = "none";
defparam \output_path_gen[0].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[0].ddio_out .power_up = "low";
defparam \output_path_gen[0].ddio_out .sync_mode = "none";
defparam \output_path_gen[0].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[0].hr_to_fr_oe (
	.datainlo(!write_oe_in[1]),
	.datainhi(!write_oe_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[0] ),
	.clk(gnd),
	.dataout(\output_path_gen[0].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[0].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[0].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[0].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[0].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[0].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[0].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[0].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[0].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[0].oe_reg .power_up = "low";

cyclonev_dqs_config \dqs_config_gen[0].dqs_config_inst (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.postamblephaseinvert(\dqsenablectrlphaseinvert[0] ),
	.dqshalfratebypass(\dqshalfratebypass[0] ),
	.enadqsenablephasetransferreg(\enadqsenablephasetransferreg[0] ),
	.dataout(\dqs_config_gen[0].dqs_config_inst~dataout ),
	.postamblephasesetting(\dqs_config_gen[0].dqs_config_inst_POSTAMBLEPHASESETTING_bus ),
	.dqsbusoutdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSBUSOUTDELAYSETTING_bus ),
	.octdelaysetting(\dqs_config_gen[0].dqs_config_inst_OCTDELAYSETTING_bus ),
	.dqsenablegatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEGATINGDELAYSETTING_bus ),
	.dqsenableungatingdelaysetting(\dqs_config_gen[0].dqs_config_inst_DQSENABLEUNGATINGDELAYSETTING_bus ));

cyclonev_ddio_out hr_to_fr_os_oct(
	.datainlo(oct_ena_in[1]),
	.datainhi(oct_ena_in[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(fr_os_oct),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oct.async_mode = "none";
defparam hr_to_fr_os_oct.half_rate_mode = "true";
defparam hr_to_fr_os_oct.power_up = "low";
defparam hr_to_fr_os_oct.sync_mode = "none";
defparam hr_to_fr_os_oct.use_new_clocking_model = "true";

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(config_clock_in),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_clk_phase_select clk_phase_select_dqs(
	.phaseinvertctrl(gnd),
	.dqsin(gnd),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(dqs_shifted_clock));
defparam clk_phase_select_dqs.invert_phase = "false";
defparam clk_phase_select_dqs.phase_setting = 0;
defparam clk_phase_select_dqs.physical_clock_source = "dqs";
defparam clk_phase_select_dqs.use_dqs_input = "false";
defparam clk_phase_select_dqs.use_phasectrlin = "false";

cyclonev_ddio_oe os_oct_ddio_oe(
	.oe(fr_os_oct),
	.clk(dqs_shifted_clock),
	.ena(vcc),
	.octreadcontrol(lfifo_oct),
	.areset(gnd),
	.sreset(gnd),
	.dataout(predelayed_os_oct),
	.dfflo(),
	.dffhi());
defparam os_oct_ddio_oe.async_mode = "none";
defparam os_oct_ddio_oe.disable_second_level_register = "true";
defparam os_oct_ddio_oe.power_up = "low";
defparam os_oct_ddio_oe.sync_mode = "none";

cyclonev_io_config \pad_gen[1].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[1] ),
	.dataout(\pad_gen[1].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[1].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[1].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[1].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[1].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[1].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_lo (
	.datainlo(write_data_in[7]),
	.datainhi(write_data_in[5]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_hi (
	.datainlo(write_data_in[6]),
	.datainhi(write_data_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].ddio_out (
	.datainlo(\output_path_gen[1].fr_data_lo ),
	.datainhi(\output_path_gen[1].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[1].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].ddio_out .async_mode = "none";
defparam \output_path_gen[1].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[1].ddio_out .power_up = "low";
defparam \output_path_gen[1].ddio_out .sync_mode = "none";
defparam \output_path_gen[1].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[1].hr_to_fr_oe (
	.datainlo(!write_oe_in[3]),
	.datainhi(!write_oe_in[2]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[1] ),
	.clk(gnd),
	.dataout(\output_path_gen[1].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[1].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[1].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[1].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[1].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[1].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[1].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[1].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[1].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[1].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[2].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[2] ),
	.dataout(\pad_gen[2].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[2].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[2].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[2].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[2].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[2].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_lo (
	.datainlo(write_data_in[11]),
	.datainhi(write_data_in[9]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_hi (
	.datainlo(write_data_in[10]),
	.datainhi(write_data_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].ddio_out (
	.datainlo(\output_path_gen[2].fr_data_lo ),
	.datainhi(\output_path_gen[2].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[2].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].ddio_out .async_mode = "none";
defparam \output_path_gen[2].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[2].ddio_out .power_up = "low";
defparam \output_path_gen[2].ddio_out .sync_mode = "none";
defparam \output_path_gen[2].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[2].hr_to_fr_oe (
	.datainlo(!write_oe_in[5]),
	.datainhi(!write_oe_in[4]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[2] ),
	.clk(gnd),
	.dataout(\output_path_gen[2].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[2].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[2].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[2].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[2].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[2].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[2].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[2].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[2].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[2].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[3].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[3] ),
	.dataout(\pad_gen[3].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[3].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[3].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[3].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[3].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[3].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_lo (
	.datainlo(write_data_in[15]),
	.datainhi(write_data_in[13]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_hi (
	.datainlo(write_data_in[14]),
	.datainhi(write_data_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].ddio_out (
	.datainlo(\output_path_gen[3].fr_data_lo ),
	.datainhi(\output_path_gen[3].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[3].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].ddio_out .async_mode = "none";
defparam \output_path_gen[3].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[3].ddio_out .power_up = "low";
defparam \output_path_gen[3].ddio_out .sync_mode = "none";
defparam \output_path_gen[3].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[3].hr_to_fr_oe (
	.datainlo(!write_oe_in[7]),
	.datainhi(!write_oe_in[6]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[3] ),
	.clk(gnd),
	.dataout(\output_path_gen[3].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[3].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[3].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[3].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[3].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[3].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[3].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[3].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[3].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[3].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[4].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[4] ),
	.dataout(\pad_gen[4].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[4].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[4].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[4].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[4].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[4].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_lo (
	.datainlo(write_data_in[19]),
	.datainhi(write_data_in[17]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_hi (
	.datainlo(write_data_in[18]),
	.datainhi(write_data_in[16]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].ddio_out (
	.datainlo(\output_path_gen[4].fr_data_lo ),
	.datainhi(\output_path_gen[4].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[4].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].ddio_out .async_mode = "none";
defparam \output_path_gen[4].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[4].ddio_out .power_up = "low";
defparam \output_path_gen[4].ddio_out .sync_mode = "none";
defparam \output_path_gen[4].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[4].hr_to_fr_oe (
	.datainlo(!write_oe_in[9]),
	.datainhi(!write_oe_in[8]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[4] ),
	.clk(gnd),
	.dataout(\output_path_gen[4].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[4].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[4].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[4].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[4].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[4].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[4].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[4].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[4].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[4].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[5].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[5] ),
	.dataout(\pad_gen[5].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[5].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[5].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[5].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[5].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[5].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_lo (
	.datainlo(write_data_in[23]),
	.datainhi(write_data_in[21]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_hi (
	.datainlo(write_data_in[22]),
	.datainhi(write_data_in[20]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].ddio_out (
	.datainlo(\output_path_gen[5].fr_data_lo ),
	.datainhi(\output_path_gen[5].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[5].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].ddio_out .async_mode = "none";
defparam \output_path_gen[5].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[5].ddio_out .power_up = "low";
defparam \output_path_gen[5].ddio_out .sync_mode = "none";
defparam \output_path_gen[5].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[5].hr_to_fr_oe (
	.datainlo(!write_oe_in[11]),
	.datainhi(!write_oe_in[10]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[5] ),
	.clk(gnd),
	.dataout(\output_path_gen[5].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[5].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[5].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[5].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[5].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[5].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[5].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[5].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[5].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[5].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[6].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[6] ),
	.dataout(\pad_gen[6].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[6].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[6].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[6].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[6].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[6].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_lo (
	.datainlo(write_data_in[27]),
	.datainhi(write_data_in[25]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_hi (
	.datainlo(write_data_in[26]),
	.datainhi(write_data_in[24]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].ddio_out (
	.datainlo(\output_path_gen[6].fr_data_lo ),
	.datainhi(\output_path_gen[6].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[6].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].ddio_out .async_mode = "none";
defparam \output_path_gen[6].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[6].ddio_out .power_up = "low";
defparam \output_path_gen[6].ddio_out .sync_mode = "none";
defparam \output_path_gen[6].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[6].hr_to_fr_oe (
	.datainlo(!write_oe_in[13]),
	.datainhi(!write_oe_in[12]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[6] ),
	.clk(gnd),
	.dataout(\output_path_gen[6].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[6].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[6].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[6].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[6].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[6].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[6].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[6].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[6].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[6].oe_reg .power_up = "low";

cyclonev_io_config \pad_gen[7].config_1 (
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(\dq_outputhalfratebypass[7] ),
	.dataout(\pad_gen[7].config_1~dataout ),
	.readfiforeadclockselect(\pad_gen[7].config_1_READFIFOREADCLOCKSELECT_bus ),
	.readfifomode(\pad_gen[7].config_1_READFIFOMODE_bus ),
	.outputregdelaysetting(\pad_gen[7].config_1_OUTPUTREGDELAYSETTING_bus ),
	.outputenabledelaysetting(\pad_gen[7].config_1_OUTPUTENABLEDELAYSETTING_bus ),
	.padtoinputregisterdelaysetting(\pad_gen[7].config_1_PADTOINPUTREGISTERDELAYSETTING_bus ));

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_lo (
	.datainlo(write_data_in[31]),
	.datainhi(write_data_in[29]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_lo ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_lo .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_lo .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_lo .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_lo .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_hi (
	.datainlo(write_data_in[30]),
	.datainhi(write_data_in[28]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_data_hi ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_hi .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_hi .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_hi .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_hi .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].ddio_out (
	.datainlo(\output_path_gen[7].fr_data_lo ),
	.datainhi(\output_path_gen[7].fr_data_hi ),
	.clkhi(dq_shifted_clock),
	.clklo(dq_shifted_clock),
	.muxsel(dq_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(\pad_gen[7].predelayed_data ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].ddio_out .async_mode = "none";
defparam \output_path_gen[7].ddio_out .half_rate_mode = "false";
defparam \output_path_gen[7].ddio_out .power_up = "low";
defparam \output_path_gen[7].ddio_out .sync_mode = "none";
defparam \output_path_gen[7].ddio_out .use_new_clocking_model = "true";

cyclonev_ddio_out \output_path_gen[7].hr_to_fr_oe (
	.datainlo(!write_oe_in[15]),
	.datainhi(!write_oe_in[14]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dq_outputhalfratebypass[7] ),
	.clk(gnd),
	.dataout(\output_path_gen[7].fr_oe ),
	.dfflo(),
	.dffhi());
defparam \output_path_gen[7].hr_to_fr_oe .async_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .half_rate_mode = "true";
defparam \output_path_gen[7].hr_to_fr_oe .power_up = "low";
defparam \output_path_gen[7].hr_to_fr_oe .sync_mode = "none";
defparam \output_path_gen[7].hr_to_fr_oe .use_new_clocking_model = "true";

dffeas \output_path_gen[7].oe_reg (
	.clk(dq_shifted_clock),
	.d(\output_path_gen[7].fr_oe ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\output_path_gen[7].oe_reg~q ),
	.prn(vcc));
defparam \output_path_gen[7].oe_reg .is_wysiwyg = "true";
defparam \output_path_gen[7].oe_reg .power_up = "low";

cyclonev_ddio_out hr_to_fr_os_lo(
	.datainlo(write_strobe[3]),
	.datainhi(write_strobe[1]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_lo),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_lo.async_mode = "none";
defparam hr_to_fr_os_lo.half_rate_mode = "true";
defparam hr_to_fr_os_lo.power_up = "low";
defparam hr_to_fr_os_lo.sync_mode = "none";
defparam hr_to_fr_os_lo.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_os_hi(
	.datainlo(write_strobe[2]),
	.datainhi(write_strobe[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_hi),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_hi.async_mode = "none";
defparam hr_to_fr_os_hi.half_rate_mode = "true";
defparam hr_to_fr_os_hi.power_up = "low";
defparam hr_to_fr_os_hi.sync_mode = "none";
defparam hr_to_fr_os_hi.use_new_clocking_model = "true";

cyclonev_ddio_out phase_align_os(
	.datainlo(fr_os_lo),
	.datainhi(fr_os_hi),
	.clkhi(dqs_shifted_clock),
	.clklo(dqs_shifted_clock),
	.muxsel(dqs_shifted_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(predelayed_os),
	.dfflo(),
	.dffhi());
defparam phase_align_os.async_mode = "none";
defparam phase_align_os.half_rate_mode = "false";
defparam phase_align_os.power_up = "low";
defparam phase_align_os.sync_mode = "none";
defparam phase_align_os.use_new_clocking_model = "true";

cyclonev_io_config dqs_io_config_1(
	.datain(gnd),
	.clk(config_clock_in),
	.ena(gnd),
	.update(gnd),
	.outputhalfratebypass(),
	.dataout(\dqs_io_config_1~dataout ),
	.readfiforeadclockselect(),
	.readfifomode(),
	.outputregdelaysetting(dqs_io_config_1_OUTPUTREGDELAYSETTING_bus),
	.outputenabledelaysetting(dqs_io_config_1_OUTPUTENABLEDELAYSETTING_bus),
	.padtoinputregisterdelaysetting());

cyclonev_delay_chain dqs_out_delay_1(
	.datain(predelayed_os),
	.delayctrlin({\dqs_outputdelaysetting_dlc[4] ,\dqs_outputdelaysetting_dlc[3] ,\dqs_outputdelaysetting_dlc[2] ,\dqs_outputdelaysetting_dlc[1] ,\dqs_outputdelaysetting_dlc[0] }),
	.dataout(os_delayed2));
defparam dqs_out_delay_1.sim_falling_delay_increment = 10;
defparam dqs_out_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_out_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_out_delay_1.sim_rising_delay_increment = 10;

cyclonev_ddio_out hr_to_fr_os_oe(
	.datainlo(!output_strobe_ena[1]),
	.datainhi(!output_strobe_ena[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(vcc),
	.clk(gnd),
	.dataout(fr_os_oe),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_os_oe.async_mode = "none";
defparam hr_to_fr_os_oe.half_rate_mode = "true";
defparam hr_to_fr_os_oe.power_up = "low";
defparam hr_to_fr_os_oe.sync_mode = "none";
defparam hr_to_fr_os_oe.use_new_clocking_model = "true";

dffeas os_oe_reg(
	.clk(dqs_shifted_clock),
	.d(fr_os_oe),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\os_oe_reg~q ),
	.prn(vcc));
defparam os_oe_reg.is_wysiwyg = "true";
defparam os_oe_reg.power_up = "low";

cyclonev_delay_chain oe_delay_1(
	.datain(\os_oe_reg~q ),
	.delayctrlin({\dqs_outputenabledelaysetting_dlc[4] ,\dqs_outputenabledelaysetting_dlc[3] ,\dqs_outputenabledelaysetting_dlc[2] ,\dqs_outputenabledelaysetting_dlc[1] ,\dqs_outputenabledelaysetting_dlc[0] }),
	.dataout(delayed_os_oe));
defparam oe_delay_1.sim_falling_delay_increment = 10;
defparam oe_delay_1.sim_intrinsic_falling_delay = 0;
defparam oe_delay_1.sim_intrinsic_rising_delay = 0;
defparam oe_delay_1.sim_rising_delay_increment = 10;

cyclonev_read_fifo_read_clock_select \input_path_gen[0].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[1] ,\rfifo_clock_select[0] }),
	.clkout(\input_path_gen[0].rfifo_rd_clk ));

cyclonev_ddio_out hr_to_fr_vfifo_inc_wr_ptr(
	.datainlo(vfifo_inc_wr_ptr[1]),
	.datainhi(vfifo_inc_wr_ptr[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_inc_wr_ptr_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_inc_wr_ptr.async_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.half_rate_mode = "true";
defparam hr_to_fr_vfifo_inc_wr_ptr.power_up = "low";
defparam hr_to_fr_vfifo_inc_wr_ptr.sync_mode = "none";
defparam hr_to_fr_vfifo_inc_wr_ptr.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_vfifo_qvld(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(vfifo_qvld_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_vfifo_qvld.async_mode = "none";
defparam hr_to_fr_vfifo_qvld.half_rate_mode = "true";
defparam hr_to_fr_vfifo_qvld.power_up = "low";
defparam hr_to_fr_vfifo_qvld.sync_mode = "none";
defparam hr_to_fr_vfifo_qvld.use_new_clocking_model = "true";

cyclonev_clk_phase_select clk_phase_select_pst_0p(
	.phaseinvertctrl(gnd),
	.dqsin(dqsbusout),
	.clkin({gnd,gnd,gnd,\leveled_dqs_clocks[0] }),
	.phasectrlin(2'b00),
	.clkout(ena_zero_phase_clock));
defparam clk_phase_select_pst_0p.invert_phase = "false";
defparam clk_phase_select_pst_0p.phase_setting = 0;
defparam clk_phase_select_pst_0p.physical_clock_source = "pst_0p";
defparam clk_phase_select_pst_0p.use_dqs_input = "false";
defparam clk_phase_select_pst_0p.use_phasectrlin = "false";

cyclonev_vfifo vfifo(
	.incwrptr(vfifo_inc_wr_ptr_fr),
	.qvldin(vfifo_qvld_fr),
	.rdclk(ena_zero_phase_clock),
	.rstn(vfifo_reset_n),
	.wrclk(dqs_shifted_clock),
	.qvldreg(dqs_pre_delayed));

cyclonev_clk_phase_select clk_phase_select_pst(
	.phaseinvertctrl(\dqsenablectrlphaseinvert[0] ),
	.dqsin(gnd),
	.clkin({\leveled_dqs_clocks[3] ,\leveled_dqs_clocks[2] ,\leveled_dqs_clocks[1] ,\leveled_dqs_clocks[0] }),
	.phasectrlin({\dqsenablectrlphasesetting[0][1] ,\dqsenablectrlphasesetting[0][0] }),
	.clkout(ena_clock));
defparam clk_phase_select_pst.invert_phase = "dynamic";
defparam clk_phase_select_pst.phase_setting = 0;
defparam clk_phase_select_pst.physical_clock_source = "pst";
defparam clk_phase_select_pst.use_dqs_input = "false";
defparam clk_phase_select_pst.use_phasectrlin = "true";

cyclonev_dqs_enable_ctrl dqs_enable_ctrl(
	.rstn(gnd),
	.dqsenablein(dqs_pre_delayed),
	.zerophaseclk(ena_zero_phase_clock),
	.enaphasetransferreg(\enadqsenablephasetransferreg[0] ),
	.levelingclk(ena_clock),
	.dqsenableout(dqs_enable_shifted));
defparam dqs_enable_ctrl.add_phase_transfer_reg = "dynamic";
defparam dqs_enable_ctrl.delay_dqs_enable = "one_and_half_cycle";

cyclonev_delay_chain dqs_ena_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsenabledelaysetting_dlc[0][4] ,\dqsenabledelaysetting_dlc[0][3] ,\dqsenabledelaysetting_dlc[0][2] ,\dqsenabledelaysetting_dlc[0][1] ,\dqsenabledelaysetting_dlc[0][0] }),
	.dataout(dqs_enable_int));
defparam dqs_ena_delay_1.sim_falling_delay_increment = 10;
defparam dqs_ena_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_ena_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_ena_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain dqs_dis_delay_1(
	.datain(dqs_enable_shifted),
	.delayctrlin({\dqsdisabledelaysetting_dlc[0][4] ,\dqsdisabledelaysetting_dlc[0][3] ,\dqsdisabledelaysetting_dlc[0][2] ,\dqsdisabledelaysetting_dlc[0][1] ,\dqsdisabledelaysetting_dlc[0][0] }),
	.dataout(dqs_disable_int));
defparam dqs_dis_delay_1.sim_falling_delay_increment = 10;
defparam dqs_dis_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_dis_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_dis_delay_1.sim_rising_delay_increment = 10;

cyclonev_dqs_delay_chain dqs_delay_chain(
	.dqsin(dqsin),
	.dqsenable(dqs_enable_int),
	.dqsdisablen(dqs_disable_int),
	.dqsupdateen(gnd),
	.testin(gnd),
	.delayctrlin({dll_delayctrl_in[6],dll_delayctrl_in[5],dll_delayctrl_in[4],dll_delayctrl_in[3],dll_delayctrl_in[2],dll_delayctrl_in[1],dll_delayctrl_in[0]}),
	.dqsbusout(dqs_shifted));
defparam dqs_delay_chain.dqs_ctrl_latches_enable = "false";
defparam dqs_delay_chain.dqs_delay_chain_bypass = "true";
defparam dqs_delay_chain.dqs_delay_chain_test_mode = "off";
defparam dqs_delay_chain.dqs_input_frequency = "0";
defparam dqs_delay_chain.dqs_phase_shift = 0;
defparam dqs_delay_chain.sim_buffer_delay_increment = 10;
defparam dqs_delay_chain.sim_buffer_intrinsic_delay = 175;

cyclonev_delay_chain dqs_in_delay_1(
	.datain(dqs_shifted),
	.delayctrlin({\dqsbusoutdelaysetting_dlc[0][4] ,\dqsbusoutdelaysetting_dlc[0][3] ,\dqsbusoutdelaysetting_dlc[0][2] ,\dqsbusoutdelaysetting_dlc[0][1] ,\dqsbusoutdelaysetting_dlc[0][0] }),
	.dataout(dqsbusout));
defparam dqs_in_delay_1.sim_falling_delay_increment = 10;
defparam dqs_in_delay_1.sim_intrinsic_falling_delay = 0;
defparam dqs_in_delay_1.sim_intrinsic_rising_delay = 0;
defparam dqs_in_delay_1.sim_rising_delay_increment = 10;

cyclonev_delay_chain \pad_gen[0].in_delay_1 (
	.datain(pad_gen0raw_input),
	.delayctrlin({\pad_gen[0].dq_inputdelaysetting_dlc[4] ,\pad_gen[0].dq_inputdelaysetting_dlc[3] ,\pad_gen[0].dq_inputdelaysetting_dlc[2] ,\pad_gen[0].dq_inputdelaysetting_dlc[1] ,\pad_gen[0].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[0] ));
defparam \pad_gen[0].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[0].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[0].capture_reg (
	.datain(\ddr_data[0] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[0].aligned_input[0] ),
	.regouthi(\input_path_gen[0].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[0].capture_reg .async_mode = "none";
defparam \input_path_gen[0].capture_reg .power_up = "low";
defparam \input_path_gen[0].capture_reg .sync_mode = "none";
defparam \input_path_gen[0].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[1].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[3] ,\rfifo_clock_select[2] }),
	.clkout(\input_path_gen[1].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[1].in_delay_1 (
	.datain(pad_gen1raw_input),
	.delayctrlin({\pad_gen[1].dq_inputdelaysetting_dlc[4] ,\pad_gen[1].dq_inputdelaysetting_dlc[3] ,\pad_gen[1].dq_inputdelaysetting_dlc[2] ,\pad_gen[1].dq_inputdelaysetting_dlc[1] ,\pad_gen[1].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[1] ));
defparam \pad_gen[1].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[1].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[1].capture_reg (
	.datain(\ddr_data[1] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[1].aligned_input[0] ),
	.regouthi(\input_path_gen[1].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[1].capture_reg .async_mode = "none";
defparam \input_path_gen[1].capture_reg .power_up = "low";
defparam \input_path_gen[1].capture_reg .sync_mode = "none";
defparam \input_path_gen[1].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[2].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[5] ,\rfifo_clock_select[4] }),
	.clkout(\input_path_gen[2].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[2].in_delay_1 (
	.datain(pad_gen2raw_input),
	.delayctrlin({\pad_gen[2].dq_inputdelaysetting_dlc[4] ,\pad_gen[2].dq_inputdelaysetting_dlc[3] ,\pad_gen[2].dq_inputdelaysetting_dlc[2] ,\pad_gen[2].dq_inputdelaysetting_dlc[1] ,\pad_gen[2].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[2] ));
defparam \pad_gen[2].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[2].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[2].capture_reg (
	.datain(\ddr_data[2] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[2].aligned_input[0] ),
	.regouthi(\input_path_gen[2].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[2].capture_reg .async_mode = "none";
defparam \input_path_gen[2].capture_reg .power_up = "low";
defparam \input_path_gen[2].capture_reg .sync_mode = "none";
defparam \input_path_gen[2].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[3].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[7] ,\rfifo_clock_select[6] }),
	.clkout(\input_path_gen[3].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[3].in_delay_1 (
	.datain(pad_gen3raw_input),
	.delayctrlin({\pad_gen[3].dq_inputdelaysetting_dlc[4] ,\pad_gen[3].dq_inputdelaysetting_dlc[3] ,\pad_gen[3].dq_inputdelaysetting_dlc[2] ,\pad_gen[3].dq_inputdelaysetting_dlc[1] ,\pad_gen[3].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[3] ));
defparam \pad_gen[3].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[3].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[3].capture_reg (
	.datain(\ddr_data[3] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[3].aligned_input[0] ),
	.regouthi(\input_path_gen[3].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[3].capture_reg .async_mode = "none";
defparam \input_path_gen[3].capture_reg .power_up = "low";
defparam \input_path_gen[3].capture_reg .sync_mode = "none";
defparam \input_path_gen[3].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[4].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[9] ,\rfifo_clock_select[8] }),
	.clkout(\input_path_gen[4].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[4].in_delay_1 (
	.datain(pad_gen4raw_input),
	.delayctrlin({\pad_gen[4].dq_inputdelaysetting_dlc[4] ,\pad_gen[4].dq_inputdelaysetting_dlc[3] ,\pad_gen[4].dq_inputdelaysetting_dlc[2] ,\pad_gen[4].dq_inputdelaysetting_dlc[1] ,\pad_gen[4].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[4] ));
defparam \pad_gen[4].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[4].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[4].capture_reg (
	.datain(\ddr_data[4] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[4].aligned_input[0] ),
	.regouthi(\input_path_gen[4].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[4].capture_reg .async_mode = "none";
defparam \input_path_gen[4].capture_reg .power_up = "low";
defparam \input_path_gen[4].capture_reg .sync_mode = "none";
defparam \input_path_gen[4].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[5].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[11] ,\rfifo_clock_select[10] }),
	.clkout(\input_path_gen[5].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[5].in_delay_1 (
	.datain(pad_gen5raw_input),
	.delayctrlin({\pad_gen[5].dq_inputdelaysetting_dlc[4] ,\pad_gen[5].dq_inputdelaysetting_dlc[3] ,\pad_gen[5].dq_inputdelaysetting_dlc[2] ,\pad_gen[5].dq_inputdelaysetting_dlc[1] ,\pad_gen[5].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[5] ));
defparam \pad_gen[5].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[5].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[5].capture_reg (
	.datain(\ddr_data[5] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[5].aligned_input[0] ),
	.regouthi(\input_path_gen[5].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[5].capture_reg .async_mode = "none";
defparam \input_path_gen[5].capture_reg .power_up = "low";
defparam \input_path_gen[5].capture_reg .sync_mode = "none";
defparam \input_path_gen[5].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[6].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[13] ,\rfifo_clock_select[12] }),
	.clkout(\input_path_gen[6].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[6].in_delay_1 (
	.datain(pad_gen6raw_input),
	.delayctrlin({\pad_gen[6].dq_inputdelaysetting_dlc[4] ,\pad_gen[6].dq_inputdelaysetting_dlc[3] ,\pad_gen[6].dq_inputdelaysetting_dlc[2] ,\pad_gen[6].dq_inputdelaysetting_dlc[1] ,\pad_gen[6].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[6] ));
defparam \pad_gen[6].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[6].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[6].capture_reg (
	.datain(\ddr_data[6] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[6].aligned_input[0] ),
	.regouthi(\input_path_gen[6].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[6].capture_reg .async_mode = "none";
defparam \input_path_gen[6].capture_reg .power_up = "low";
defparam \input_path_gen[6].capture_reg .sync_mode = "none";
defparam \input_path_gen[6].capture_reg .use_clkn = "false";

cyclonev_read_fifo_read_clock_select \input_path_gen[7].read_fifo_clk_sel (
	.clkin({hr_seq_clock,dqs_shifted_clock,GND_port}),
	.clksel({\rfifo_clock_select[15] ,\rfifo_clock_select[14] }),
	.clkout(\input_path_gen[7].rfifo_rd_clk ));

cyclonev_delay_chain \pad_gen[7].in_delay_1 (
	.datain(pad_gen7raw_input),
	.delayctrlin({\pad_gen[7].dq_inputdelaysetting_dlc[4] ,\pad_gen[7].dq_inputdelaysetting_dlc[3] ,\pad_gen[7].dq_inputdelaysetting_dlc[2] ,\pad_gen[7].dq_inputdelaysetting_dlc[1] ,\pad_gen[7].dq_inputdelaysetting_dlc[0] }),
	.dataout(\ddr_data[7] ));
defparam \pad_gen[7].in_delay_1 .sim_falling_delay_increment = 10;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_falling_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_intrinsic_rising_delay = 200;
defparam \pad_gen[7].in_delay_1 .sim_rising_delay_increment = 10;

cyclonev_ddio_in \input_path_gen[7].capture_reg (
	.datain(\ddr_data[7] ),
	.clk(!dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(\input_path_gen[7].aligned_input[0] ),
	.regouthi(\input_path_gen[7].aligned_input[1] ),
	.dfflo());
defparam \input_path_gen[7].capture_reg .async_mode = "none";
defparam \input_path_gen[7].capture_reg .power_up = "low";
defparam \input_path_gen[7].capture_reg .sync_mode = "none";
defparam \input_path_gen[7].capture_reg .use_clkn = "false";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en(
	.datainlo(lfifo_rdata_en[1]),
	.datainhi(lfifo_rdata_en[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en.use_new_clocking_model = "true";

cyclonev_ddio_out hr_to_fr_lfifo_rdata_en_full(
	.datainlo(lfifo_rdata_en_full[1]),
	.datainhi(lfifo_rdata_en_full[0]),
	.clkhi(hr_seq_clock),
	.clklo(hr_seq_clock),
	.muxsel(hr_seq_clock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.hrbypass(\dqshalfratebypass[0] ),
	.clk(gnd),
	.dataout(lfifo_rdata_en_full_fr),
	.dfflo(),
	.dffhi());
defparam hr_to_fr_lfifo_rdata_en_full.async_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.half_rate_mode = "true";
defparam hr_to_fr_lfifo_rdata_en_full.power_up = "low";
defparam hr_to_fr_lfifo_rdata_en_full.sync_mode = "none";
defparam hr_to_fr_lfifo_rdata_en_full.use_new_clocking_model = "true";

endmodule

module terminal_qsys_hps_sdram_p0_acv_ldc_25 (
	pll_dqs_clk,
	pll_hr_clk,
	afi_clk,
	avl_clk,
	dll_phy_delayctrl)/* synthesis synthesis_greybox=0 */;
input 	pll_dqs_clk;
input 	pll_hr_clk;
output 	afi_clk;
output 	avl_clk;
input 	[6:0] dll_phy_delayctrl;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \leveled_dqs_clocks[1] ;
wire \leveled_dqs_clocks[2] ;
wire \leveled_dqs_clocks[3] ;
wire \leveled_hr_clocks[1] ;
wire \leveled_hr_clocks[2] ;
wire \leveled_hr_clocks[3] ;

wire [3:0] leveling_delay_chain_dqs_CLKOUT_bus;
wire [3:0] leveling_delay_chain_hr_CLKOUT_bus;

assign afi_clk = leveling_delay_chain_dqs_CLKOUT_bus[0];
assign \leveled_dqs_clocks[1]  = leveling_delay_chain_dqs_CLKOUT_bus[1];
assign \leveled_dqs_clocks[2]  = leveling_delay_chain_dqs_CLKOUT_bus[2];
assign \leveled_dqs_clocks[3]  = leveling_delay_chain_dqs_CLKOUT_bus[3];

assign avl_clk = leveling_delay_chain_hr_CLKOUT_bus[0];
assign \leveled_hr_clocks[1]  = leveling_delay_chain_hr_CLKOUT_bus[1];
assign \leveled_hr_clocks[2]  = leveling_delay_chain_hr_CLKOUT_bus[2];
assign \leveled_hr_clocks[3]  = leveling_delay_chain_hr_CLKOUT_bus[3];

cyclonev_leveling_delay_chain leveling_delay_chain_dqs(
	.clkin(pll_dqs_clk),
	.delayctrlin({dll_phy_delayctrl[6],dll_phy_delayctrl[5],dll_phy_delayctrl[4],dll_phy_delayctrl[3],dll_phy_delayctrl[2],dll_phy_delayctrl[1],dll_phy_delayctrl[0]}),
	.clkout(leveling_delay_chain_dqs_CLKOUT_bus));
defparam leveling_delay_chain_dqs.physical_clock_source = "dqs";
defparam leveling_delay_chain_dqs.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_dqs.sim_buffer_intrinsic_delay = 175;

cyclonev_leveling_delay_chain leveling_delay_chain_hr(
	.clkin(pll_dqs_clk),
	.delayctrlin(7'b0000000),
	.clkout(leveling_delay_chain_hr_CLKOUT_bus));
defparam leveling_delay_chain_hr.physical_clock_source = "hr";
defparam leveling_delay_chain_hr.sim_buffer_delay_increment = 10;
defparam leveling_delay_chain_hr.sim_buffer_intrinsic_delay = 175;

endmodule

module terminal_qsys_hps_sdram_pll (
	pll_mem_clk,
	pll_write_clk)/* synthesis synthesis_greybox=0 */;
output 	pll_mem_clk;
output 	pll_write_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_out[2] ;
wire \clk_out[3] ;

wire [3:0] pll_CLK_OUT_bus;

assign pll_mem_clk = pll_CLK_OUT_bus[0];
assign pll_write_clk = pll_CLK_OUT_bus[1];
assign \clk_out[2]  = pll_CLK_OUT_bus[2];
assign \clk_out[3]  = pll_CLK_OUT_bus[3];

cyclonev_hps_sdram_pll pll(
	.ref_clk(gnd),
	.clk_out(pll_CLK_OUT_bus));

endmodule

module terminal_qsys_terminal_qsys_leds (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	wait_latency_counter_1,
	wait_latency_counter_0,
	reset_n,
	writedata,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	clk)/* synthesis synthesis_greybox=0 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	reset_n;
input 	[31:0] writedata;
input 	m0_write;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'h4040404040404040;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'h4040404040404040;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'h4040404040404040;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'h4040404040404040;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'h4040404040404040;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'h4040404040404040;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'h4040404040404040;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'h4040404040404040;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \readdata[8] (
	.dataa(!data_out_8),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[8] .extended_lut = "off";
defparam \readdata[8] .lut_mask = 64'h4040404040404040;
defparam \readdata[8] .shared_arith = "off";

cyclonev_lcell_comb \readdata[9] (
	.dataa(!data_out_9),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[9] .extended_lut = "off";
defparam \readdata[9] .lut_mask = 64'h4040404040404040;
defparam \readdata[9] .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(!int_nxt_addr_reg_dly_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h0800000008000000;
defparam \always0~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0 (
	h2f_lw_ARVALID_0,
	h2f_lw_AWVALID_0,
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARADDR_15,
	h2f_lw_ARADDR_16,
	h2f_lw_ARADDR_17,
	h2f_lw_ARADDR_18,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWADDR_15,
	h2f_lw_AWADDR_16,
	h2f_lw_AWADDR_17,
	h2f_lw_AWADDR_18,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	wait_latency_counter_1,
	wait_latency_counter_0,
	wait_latency_counter_11,
	wait_latency_counter_01,
	wait_latency_counter_12,
	wait_latency_counter_02,
	cmd_sink_ready,
	nonposted_cmd_accepted,
	WideOr1,
	src_payload_0,
	WideOr11,
	nonposted_cmd_accepted1,
	src_payload,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_data_0,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_6,
	src_data_7,
	src_data_8,
	src_data_9,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	src_payload33,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	in_data_reg_0,
	altera_reset_synchronizer_int_chain_out,
	m0_write,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	in_data_reg_01,
	altera_reset_synchronizer_int_chain_out1,
	m0_write1,
	int_nxt_addr_reg_dly_31,
	int_nxt_addr_reg_dly_21,
	in_data_reg_110,
	in_data_reg_210,
	in_data_reg_32,
	in_data_reg_41,
	in_data_reg_51,
	in_data_reg_61,
	in_data_reg_71,
	in_data_reg_81,
	in_data_reg_91,
	in_data_reg_101,
	in_data_reg_111,
	in_data_reg_121,
	in_data_reg_131,
	in_data_reg_141,
	in_data_reg_151,
	in_data_reg_161,
	in_data_reg_171,
	in_data_reg_181,
	in_data_reg_191,
	in_data_reg_201,
	in_data_reg_211,
	in_data_reg_221,
	in_data_reg_231,
	in_data_reg_241,
	in_data_reg_251,
	in_data_reg_261,
	in_data_reg_271,
	in_data_reg_281,
	in_data_reg_291,
	in_data_reg_301,
	in_data_reg_311,
	in_data_reg_02,
	m0_write2,
	int_nxt_addr_reg_dly_32,
	int_nxt_addr_reg_dly_22,
	in_data_reg_112,
	in_data_reg_212,
	in_data_reg_33,
	in_data_reg_42,
	in_data_reg_52,
	in_data_reg_62,
	in_data_reg_72,
	in_data_reg_82,
	in_data_reg_92,
	altera_reset_synchronizer_int_chain_out2,
	readdata_0,
	readdata_01,
	readdata_02,
	readdata_03,
	readdata_04,
	readdata_1,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_2,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_3,
	readdata_31,
	readdata_32,
	readdata_33,
	readdata_34,
	readdata_4,
	readdata_41,
	readdata_42,
	readdata_43,
	readdata_44,
	readdata_5,
	readdata_51,
	readdata_52,
	readdata_53,
	readdata_54,
	readdata_6,
	readdata_61,
	readdata_62,
	readdata_63,
	readdata_64,
	readdata_7,
	readdata_71,
	readdata_72,
	readdata_73,
	readdata_74,
	readdata_8,
	readdata_81,
	readdata_82,
	readdata_83,
	readdata_84,
	readdata_9,
	readdata_91,
	readdata_92,
	readdata_93,
	readdata_94,
	readdata_10,
	readdata_101,
	readdata_102,
	readdata_111,
	readdata_112,
	readdata_113,
	readdata_121,
	readdata_122,
	readdata_123,
	readdata_131,
	readdata_132,
	readdata_133,
	readdata_141,
	readdata_142,
	readdata_143,
	readdata_15,
	readdata_151,
	readdata_152,
	readdata_16,
	readdata_161,
	readdata_162,
	readdata_17,
	readdata_171,
	readdata_172,
	readdata_18,
	readdata_181,
	readdata_182,
	readdata_19,
	readdata_191,
	readdata_192,
	readdata_20,
	readdata_201,
	readdata_202,
	readdata_211,
	readdata_212,
	readdata_213,
	readdata_221,
	readdata_222,
	readdata_223,
	readdata_231,
	readdata_232,
	readdata_233,
	readdata_241,
	readdata_242,
	readdata_243,
	readdata_25,
	readdata_251,
	readdata_252,
	readdata_26,
	readdata_261,
	readdata_262,
	readdata_27,
	readdata_271,
	readdata_272,
	readdata_28,
	readdata_281,
	readdata_282,
	readdata_29,
	readdata_291,
	readdata_292,
	readdata_30,
	readdata_301,
	readdata_302,
	readdata_311,
	readdata_312,
	readdata_313,
	int_nxt_addr_reg_dly_33,
	int_nxt_addr_reg_dly_23,
	int_nxt_addr_reg_dly_34,
	int_nxt_addr_reg_dly_24,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARADDR_5;
input 	h2f_lw_ARADDR_6;
input 	h2f_lw_ARADDR_7;
input 	h2f_lw_ARADDR_8;
input 	h2f_lw_ARADDR_9;
input 	h2f_lw_ARADDR_10;
input 	h2f_lw_ARADDR_11;
input 	h2f_lw_ARADDR_12;
input 	h2f_lw_ARADDR_13;
input 	h2f_lw_ARADDR_14;
input 	h2f_lw_ARADDR_15;
input 	h2f_lw_ARADDR_16;
input 	h2f_lw_ARADDR_17;
input 	h2f_lw_ARADDR_18;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWADDR_15;
input 	h2f_lw_AWADDR_16;
input 	h2f_lw_AWADDR_17;
input 	h2f_lw_AWADDR_18;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
output 	wait_latency_counter_12;
output 	wait_latency_counter_02;
output 	cmd_sink_ready;
output 	nonposted_cmd_accepted;
output 	WideOr1;
output 	src_payload_0;
output 	WideOr11;
output 	nonposted_cmd_accepted1;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_data_0;
output 	src_data_1;
output 	src_data_2;
output 	src_data_3;
output 	src_data_4;
output 	src_data_5;
output 	src_data_6;
output 	src_data_7;
output 	src_data_8;
output 	src_data_9;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_100;
output 	src_data_101;
output 	src_data_102;
output 	src_data_103;
output 	in_data_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
output 	in_data_reg_01;
input 	altera_reset_synchronizer_int_chain_out1;
output 	m0_write1;
output 	int_nxt_addr_reg_dly_31;
output 	int_nxt_addr_reg_dly_21;
output 	in_data_reg_110;
output 	in_data_reg_210;
output 	in_data_reg_32;
output 	in_data_reg_41;
output 	in_data_reg_51;
output 	in_data_reg_61;
output 	in_data_reg_71;
output 	in_data_reg_81;
output 	in_data_reg_91;
output 	in_data_reg_101;
output 	in_data_reg_111;
output 	in_data_reg_121;
output 	in_data_reg_131;
output 	in_data_reg_141;
output 	in_data_reg_151;
output 	in_data_reg_161;
output 	in_data_reg_171;
output 	in_data_reg_181;
output 	in_data_reg_191;
output 	in_data_reg_201;
output 	in_data_reg_211;
output 	in_data_reg_221;
output 	in_data_reg_231;
output 	in_data_reg_241;
output 	in_data_reg_251;
output 	in_data_reg_261;
output 	in_data_reg_271;
output 	in_data_reg_281;
output 	in_data_reg_291;
output 	in_data_reg_301;
output 	in_data_reg_311;
output 	in_data_reg_02;
output 	m0_write2;
output 	int_nxt_addr_reg_dly_32;
output 	int_nxt_addr_reg_dly_22;
output 	in_data_reg_112;
output 	in_data_reg_212;
output 	in_data_reg_33;
output 	in_data_reg_42;
output 	in_data_reg_52;
output 	in_data_reg_62;
output 	in_data_reg_72;
output 	in_data_reg_82;
output 	in_data_reg_92;
input 	altera_reset_synchronizer_int_chain_out2;
input 	readdata_0;
input 	readdata_01;
input 	readdata_02;
input 	readdata_03;
input 	readdata_04;
input 	readdata_1;
input 	readdata_11;
input 	readdata_12;
input 	readdata_13;
input 	readdata_14;
input 	readdata_2;
input 	readdata_21;
input 	readdata_22;
input 	readdata_23;
input 	readdata_24;
input 	readdata_3;
input 	readdata_31;
input 	readdata_32;
input 	readdata_33;
input 	readdata_34;
input 	readdata_4;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
input 	readdata_44;
input 	readdata_5;
input 	readdata_51;
input 	readdata_52;
input 	readdata_53;
input 	readdata_54;
input 	readdata_6;
input 	readdata_61;
input 	readdata_62;
input 	readdata_63;
input 	readdata_64;
input 	readdata_7;
input 	readdata_71;
input 	readdata_72;
input 	readdata_73;
input 	readdata_74;
input 	readdata_8;
input 	readdata_81;
input 	readdata_82;
input 	readdata_83;
input 	readdata_84;
input 	readdata_9;
input 	readdata_91;
input 	readdata_92;
input 	readdata_93;
input 	readdata_94;
input 	readdata_10;
input 	readdata_101;
input 	readdata_102;
input 	readdata_111;
input 	readdata_112;
input 	readdata_113;
input 	readdata_121;
input 	readdata_122;
input 	readdata_123;
input 	readdata_131;
input 	readdata_132;
input 	readdata_133;
input 	readdata_141;
input 	readdata_142;
input 	readdata_143;
input 	readdata_15;
input 	readdata_151;
input 	readdata_152;
input 	readdata_16;
input 	readdata_161;
input 	readdata_162;
input 	readdata_17;
input 	readdata_171;
input 	readdata_172;
input 	readdata_18;
input 	readdata_181;
input 	readdata_182;
input 	readdata_19;
input 	readdata_191;
input 	readdata_192;
input 	readdata_20;
input 	readdata_201;
input 	readdata_202;
input 	readdata_211;
input 	readdata_212;
input 	readdata_213;
input 	readdata_221;
input 	readdata_222;
input 	readdata_223;
input 	readdata_231;
input 	readdata_232;
input 	readdata_233;
input 	readdata_241;
input 	readdata_242;
input 	readdata_243;
input 	readdata_25;
input 	readdata_251;
input 	readdata_252;
input 	readdata_26;
input 	readdata_261;
input 	readdata_262;
input 	readdata_27;
input 	readdata_271;
input 	readdata_272;
input 	readdata_28;
input 	readdata_281;
input 	readdata_282;
input 	readdata_29;
input 	readdata_291;
input 	readdata_292;
input 	readdata_30;
input 	readdata_301;
input 	readdata_302;
input 	readdata_311;
input 	readdata_312;
input 	readdata_313;
output 	int_nxt_addr_reg_dly_33;
output 	int_nxt_addr_reg_dly_23;
output 	int_nxt_addr_reg_dly_34;
output 	int_nxt_addr_reg_dly_24;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[7]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[6]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[9]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[8]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[11]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[10]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[15]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[14]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[13]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[12]~q ;
wire \hps_h2f_lw_axi_master_agent|Add5~9_sumout ;
wire \hps_h2f_lw_axi_master_agent|Add5~13_sumout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \router_001|Equal1~0_combout ;
wire \router_001|Equal1~1_combout ;
wire \router_001|Equal5~0_combout ;
wire \cmd_mux_005|saved_grant[1]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \switches_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \switches_s1_translator|wait_latency_counter[1]~q ;
wire \switches_s1_translator|wait_latency_counter[0]~q ;
wire \switches_s1_agent|cp_ready~0_combout ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_demux_001|sink_ready~0_combout ;
wire \hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ;
wire \router_001|src_channel[4]~0_combout ;
wire \cmd_mux_003|saved_grant[1]~q ;
wire \router_001|Equal4~0_combout ;
wire \router_001|Equal4~1_combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \base_address_ddr_s1_agent|WideOr0~0_combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \base_address_ddr_s1_agent|local_write~combout ;
wire \base_address_ddr_s1_agent_rsp_fifo|write~0_combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \cmd_demux_001|sink_ready~1_combout ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \rbf_id_control_slave_translator|wait_latency_counter[1]~q ;
wire \rbf_id_control_slave_translator|wait_latency_counter[0]~q ;
wire \rbf_id_control_slave_agent|cp_ready~0_combout ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_mux|saved_grant[1]~q ;
wire \router_001|Equal1~2_combout ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \state_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \state_s1_translator|wait_latency_counter[1]~q ;
wire \state_s1_translator|wait_latency_counter[0]~q ;
wire \state_s1_agent|cp_ready~0_combout ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_mux_001|saved_grant[1]~q ;
wire \cmd_demux_001|WideOr0~0_combout ;
wire \cmd_mux_002|saved_grant[1]~q ;
wire \router_001|Equal3~0_combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \control_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \control_s1_agent|WideOr0~0_combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \control_s1_agent|local_write~combout ;
wire \control_s1_agent_rsp_fifo|write~0_combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_demux_001|sink_ready~4_combout ;
wire \cmd_mux_004|saved_grant[1]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ;
wire \leds_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ;
wire \leds_s1_agent|WideOr0~0_combout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ;
wire \leds_s1_agent|local_write~combout ;
wire \leds_s1_agent_rsp_fifo|write~0_combout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ;
wire \router_001|src_channel[4]~1_combout ;
wire \cmd_demux_001|sink_ready~5_combout ;
wire \hps_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ;
wire \hps_h2f_lw_axi_master_agent|sop_enable~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[4]~q ;
wire \router|Equal3~6_combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[18]~0_combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[17]~1_combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[16]~2_combout ;
wire \router|Equal3~7_combout ;
wire \router|Equal4~0_combout ;
wire \hps_h2f_lw_axi_master_wr_limiter|has_pending_responses~q ;
wire \hps_h2f_lw_axi_master_wr_limiter|last_channel[2]~q ;
wire \hps_h2f_lw_axi_master_wr_limiter|last_channel[4]~q ;
wire \cmd_mux_003|saved_grant[0]~q ;
wire \cmd_demux|sink_ready~0_combout ;
wire \cmd_mux_002|saved_grant[0]~q ;
wire \cmd_demux|sink_ready~1_combout ;
wire \cmd_mux_004|saved_grant[0]~q ;
wire \cmd_demux|sink_ready~2_combout ;
wire \control_s1_translator|read_latency_shift_reg[0]~q ;
wire \control_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \control_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][59]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \rsp_demux_002|src0_valid~combout ;
wire \base_address_ddr_s1_translator|read_latency_shift_reg[0]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][59]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \rsp_demux_003|src0_valid~combout ;
wire \leds_s1_translator|read_latency_shift_reg[0]~q ;
wire \leds_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][116]~q ;
wire \leds_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][59]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \rsp_demux_004|src0_valid~combout ;
wire \control_s1_agent|comb~0_combout ;
wire \rsp_demux_002|src1_valid~0_combout ;
wire \control_s1_agent_rsp_fifo|mem[0][117]~q ;
wire \control_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \control_s1_agent_rsp_fifo|mem[0][69]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][65]~q ;
wire \control_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \base_address_ddr_s1_agent|comb~0_combout ;
wire \rsp_demux_003|src1_valid~0_combout ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][117]~q ;
wire \base_address_ddr_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][69]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][65]~q ;
wire \base_address_ddr_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \leds_s1_agent|comb~0_combout ;
wire \rsp_demux_004|src1_valid~0_combout ;
wire \leds_s1_agent_rsp_fifo|mem[0][117]~q ;
wire \leds_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \leds_s1_agent_rsp_fifo|mem[0][69]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][65]~q ;
wire \leds_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \switches_s1_agent_rsp_fifo|mem[0][117]~q ;
wire \switches_s1_translator|read_latency_shift_reg[0]~q ;
wire \switches_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \switches_s1_agent_rdata_fifo|empty~combout ;
wire \switches_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \switches_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \switches_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \switches_s1_agent_rsp_fifo|mem[0][69]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][65]~q ;
wire \switches_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \state_s1_agent_rsp_fifo|mem[0][117]~q ;
wire \state_s1_translator|read_latency_shift_reg[0]~q ;
wire \state_s1_agent_rdata_fifo|mem_used[0]~q ;
wire \state_s1_agent_rdata_fifo|empty~combout ;
wire \state_s1_agent_rsp_fifo|mem[0][57]~q ;
wire \state_s1_agent_rsp_fifo|mem_used[0]~q ;
wire \state_s1_agent|uncompressor|last_packet_beat~0_combout ;
wire \state_s1_agent_rsp_fifo|mem[0][69]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][68]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][67]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][66]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][65]~q ;
wire \state_s1_agent|uncompressor|last_packet_beat~1_combout ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][117]~q ;
wire \rbf_id_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \rbf_id_control_slave_agent_rdata_fifo|mem_used[0]~q ;
wire \rbf_id_control_slave_agent_rdata_fifo|empty~combout ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][57]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem_used[0]~q ;
wire \rbf_id_control_slave_agent|uncompressor|last_packet_beat~0_combout ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][69]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][68]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][67]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][66]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][65]~q ;
wire \rbf_id_control_slave_agent|uncompressor|last_packet_beat~1_combout ;
wire \control_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][96]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][96]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][96]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][97]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][97]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][97]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][98]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][98]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][98]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][99]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][99]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][99]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][100]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][100]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][100]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][101]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][101]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][101]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][102]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][102]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][102]~q ;
wire \control_s1_agent_rsp_fifo|mem[0][103]~q ;
wire \base_address_ddr_s1_agent_rsp_fifo|mem[0][103]~q ;
wire \leds_s1_agent_rsp_fifo|mem[0][103]~q ;
wire \control_s1_translator|av_readdata_pre[0]~q ;
wire \control_s1_agent_rdata_fifo|always4~0_combout ;
wire \control_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[0]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|always4~0_combout ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \leds_s1_translator|av_readdata_pre[0]~q ;
wire \leds_s1_agent_rdata_fifo|always4~0_combout ;
wire \leds_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \state_s1_translator|av_readdata_pre[0]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][0]~q ;
wire \switches_s1_translator|av_readdata_pre[0]~q ;
wire \control_s1_translator|av_readdata_pre[1]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[1]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \leds_s1_translator|av_readdata_pre[1]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \state_s1_translator|av_readdata_pre[1]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][1]~q ;
wire \switches_s1_translator|av_readdata_pre[1]~q ;
wire \control_s1_translator|av_readdata_pre[2]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[2]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \leds_s1_translator|av_readdata_pre[2]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \state_s1_translator|av_readdata_pre[2]~q ;
wire \rbf_id_control_slave_agent_rdata_fifo|mem[0][11]~q ;
wire \rbf_id_control_slave_translator|av_readdata_pre[30]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][2]~q ;
wire \switches_s1_translator|av_readdata_pre[2]~q ;
wire \control_s1_translator|av_readdata_pre[3]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[3]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \leds_s1_translator|av_readdata_pre[3]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \state_s1_translator|av_readdata_pre[3]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][3]~q ;
wire \switches_s1_translator|av_readdata_pre[3]~q ;
wire \control_s1_translator|av_readdata_pre[4]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[4]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \leds_s1_translator|av_readdata_pre[4]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \state_s1_translator|av_readdata_pre[4]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][4]~q ;
wire \switches_s1_translator|av_readdata_pre[4]~q ;
wire \control_s1_translator|av_readdata_pre[5]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[5]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \leds_s1_translator|av_readdata_pre[5]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \state_s1_translator|av_readdata_pre[5]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][5]~q ;
wire \switches_s1_translator|av_readdata_pre[5]~q ;
wire \control_s1_translator|av_readdata_pre[6]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[6]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \leds_s1_translator|av_readdata_pre[6]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \state_s1_translator|av_readdata_pre[6]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][6]~q ;
wire \switches_s1_translator|av_readdata_pre[6]~q ;
wire \control_s1_translator|av_readdata_pre[7]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[7]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \leds_s1_translator|av_readdata_pre[7]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \state_s1_translator|av_readdata_pre[7]~q ;
wire \rbf_id_control_slave_agent_rdata_fifo|mem[0][10]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][7]~q ;
wire \switches_s1_translator|av_readdata_pre[7]~q ;
wire \control_s1_translator|av_readdata_pre[8]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[8]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \leds_s1_translator|av_readdata_pre[8]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \state_s1_translator|av_readdata_pre[8]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][8]~q ;
wire \switches_s1_translator|av_readdata_pre[8]~q ;
wire \state_s1_translator|av_readdata_pre[9]~q ;
wire \control_s1_translator|av_readdata_pre[9]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[9]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \leds_s1_translator|av_readdata_pre[9]~q ;
wire \leds_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \switches_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \switches_s1_translator|av_readdata_pre[9]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][9]~q ;
wire \control_s1_translator|av_readdata_pre[10]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][10]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[10]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][10]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][10]~q ;
wire \state_s1_translator|av_readdata_pre[10]~q ;
wire \control_s1_translator|av_readdata_pre[11]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][11]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[11]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][11]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][11]~q ;
wire \state_s1_translator|av_readdata_pre[11]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[12]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][12]~q ;
wire \control_s1_translator|av_readdata_pre[12]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][12]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][12]~q ;
wire \state_s1_translator|av_readdata_pre[12]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[13]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][13]~q ;
wire \control_s1_translator|av_readdata_pre[13]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][13]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][13]~q ;
wire \state_s1_translator|av_readdata_pre[13]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[14]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][14]~q ;
wire \control_s1_translator|av_readdata_pre[14]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][14]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][14]~q ;
wire \state_s1_translator|av_readdata_pre[14]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[15]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][15]~q ;
wire \control_s1_translator|av_readdata_pre[15]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][15]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][15]~q ;
wire \state_s1_translator|av_readdata_pre[15]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[16]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][16]~q ;
wire \control_s1_translator|av_readdata_pre[16]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][16]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][16]~q ;
wire \state_s1_translator|av_readdata_pre[16]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[17]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][17]~q ;
wire \control_s1_translator|av_readdata_pre[17]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][17]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][17]~q ;
wire \state_s1_translator|av_readdata_pre[17]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[18]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][18]~q ;
wire \control_s1_translator|av_readdata_pre[18]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][18]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][18]~q ;
wire \state_s1_translator|av_readdata_pre[18]~q ;
wire \control_s1_translator|av_readdata_pre[19]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][19]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[19]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][19]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][19]~q ;
wire \state_s1_translator|av_readdata_pre[19]~q ;
wire \control_s1_translator|av_readdata_pre[20]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][20]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[20]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][20]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][20]~q ;
wire \state_s1_translator|av_readdata_pre[20]~q ;
wire \control_s1_translator|av_readdata_pre[21]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][21]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[21]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][21]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][21]~q ;
wire \state_s1_translator|av_readdata_pre[21]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[22]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][22]~q ;
wire \control_s1_translator|av_readdata_pre[22]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][22]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][22]~q ;
wire \state_s1_translator|av_readdata_pre[22]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[23]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][23]~q ;
wire \control_s1_translator|av_readdata_pre[23]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][23]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][23]~q ;
wire \state_s1_translator|av_readdata_pre[23]~q ;
wire \control_s1_translator|av_readdata_pre[24]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][24]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[24]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][24]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][24]~q ;
wire \state_s1_translator|av_readdata_pre[24]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[25]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][25]~q ;
wire \control_s1_translator|av_readdata_pre[25]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][25]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][25]~q ;
wire \state_s1_translator|av_readdata_pre[25]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[26]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][26]~q ;
wire \control_s1_translator|av_readdata_pre[26]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][26]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][26]~q ;
wire \state_s1_translator|av_readdata_pre[26]~q ;
wire \control_s1_translator|av_readdata_pre[27]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][27]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[27]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][27]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][27]~q ;
wire \state_s1_translator|av_readdata_pre[27]~q ;
wire \control_s1_translator|av_readdata_pre[28]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][28]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[28]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][28]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][28]~q ;
wire \state_s1_translator|av_readdata_pre[28]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[29]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][29]~q ;
wire \control_s1_translator|av_readdata_pre[29]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][29]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][29]~q ;
wire \state_s1_translator|av_readdata_pre[29]~q ;
wire \control_s1_translator|av_readdata_pre[30]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][30]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[30]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][30]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][30]~q ;
wire \state_s1_translator|av_readdata_pre[30]~q ;
wire \base_address_ddr_s1_translator|av_readdata_pre[31]~q ;
wire \base_address_ddr_s1_agent_rdata_fifo|mem[0][31]~q ;
wire \control_s1_translator|av_readdata_pre[31]~q ;
wire \control_s1_agent_rdata_fifo|mem[0][31]~q ;
wire \state_s1_agent_rdata_fifo|mem[0][31]~q ;
wire \state_s1_translator|av_readdata_pre[31]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][92]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][92]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][93]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][93]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][94]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][94]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][95]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][95]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][96]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][96]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][96]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][97]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][97]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][97]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][98]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][98]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][98]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][99]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][99]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][99]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][100]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][100]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][100]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][101]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][101]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][101]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][102]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][102]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][102]~q ;
wire \switches_s1_agent_rsp_fifo|mem[0][103]~q ;
wire \rbf_id_control_slave_agent_rsp_fifo|mem[0][103]~q ;
wire \state_s1_agent_rsp_fifo|mem[0][103]~q ;
wire \hps_h2f_lw_axi_master_rd_limiter|last_channel[5]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \cmd_mux_005|last_cycle~0_combout ;
wire \switches_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \switches_s1_agent_rdata_fifo|read~0_combout ;
wire \switches_s1_agent_rsp_fifo|write~0_combout ;
wire \switches_s1_agent_rsp_fifo|write~1_combout ;
wire \hps_h2f_lw_axi_master_agent|Decoder1~0_combout ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \hps_h2f_lw_axi_master_agent|Add2~0_combout ;
wire \hps_h2f_lw_axi_master_agent|Add2~1_combout ;
wire \hps_h2f_lw_axi_master_agent|Add2~2_combout ;
wire \switches_s1_agent|cp_ready~1_combout ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_demux_001|WideOr0~combout ;
wire \router_001|src_data[90]~0_combout ;
wire \router_001|src_data[91]~1_combout ;
wire \hps_h2f_lw_axi_master_wr_limiter|last_channel[3]~q ;
wire \cmd_demux|src3_valid~0_combout ;
wire \hps_h2f_lw_axi_master_rd_limiter|last_channel[3]~q ;
wire \cmd_demux_001|src3_valid~0_combout ;
wire \cmd_demux_001|src3_valid~1_combout ;
wire \cmd_mux_003|src_valid~0_combout ;
wire \cmd_mux_003|src_payload[0]~combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \base_address_ddr_s1_agent|cp_ready~2_combout ;
wire \base_address_ddr_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \rsp_demux_003|WideOr0~0_combout ;
wire \base_address_ddr_s1_agent_rsp_fifo|read~0_combout ;
wire \cmd_mux_003|src_data[78]~combout ;
wire \cmd_mux_003|src_data[79]~combout ;
wire \cmd_mux_003|src_data[35]~combout ;
wire \cmd_mux_003|src_data[34]~combout ;
wire \cmd_mux_003|src_data[33]~combout ;
wire \cmd_mux_003|src_data[32]~combout ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ;
wire \hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ;
wire \hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ;
wire \hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ;
wire \hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ;
wire \hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ;
wire \hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ;
wire \hps_h2f_lw_axi_master_agent|write_cp_data[66]~3_combout ;
wire \hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ;
wire \hps_h2f_lw_axi_master_agent|write_cp_data[65]~4_combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \router_001|Equal1~3_combout ;
wire \hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ;
wire \rbf_id_control_slave_agent|uncompressor|last_packet_beat~2_combout ;
wire \rbf_id_control_slave_agent_rdata_fifo|read~0_combout ;
wire \rbf_id_control_slave_agent_rsp_fifo|write~0_combout ;
wire \rbf_id_control_slave_agent_rsp_fifo|write~1_combout ;
wire \cmd_mux|src_valid~0_combout ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \rbf_id_control_slave_agent|cp_ready~1_combout ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \router_001|Equal2~0_combout ;
wire \hps_h2f_lw_axi_master_rd_limiter|last_channel[1]~q ;
wire \cmd_mux_001|src_valid~0_combout ;
wire \state_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \state_s1_agent_rdata_fifo|read~0_combout ;
wire \state_s1_agent_rsp_fifo|write~0_combout ;
wire \state_s1_agent_rsp_fifo|write~1_combout ;
wire \cmd_mux_001|src_valid~1_combout ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \state_s1_agent|cp_ready~1_combout ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_demux|src2_valid~0_combout ;
wire \hps_h2f_lw_axi_master_rd_limiter|last_channel[2]~q ;
wire \cmd_demux_001|src2_valid~0_combout ;
wire \cmd_demux_001|src2_valid~1_combout ;
wire \cmd_mux_002|src_valid~0_combout ;
wire \cmd_mux_002|src_payload[0]~combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \control_s1_agent|cp_ready~2_combout ;
wire \control_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \rsp_demux_002|WideOr0~0_combout ;
wire \control_s1_agent_rsp_fifo|read~0_combout ;
wire \cmd_mux_002|src_data[78]~combout ;
wire \cmd_mux_002|src_data[79]~combout ;
wire \cmd_mux_002|src_data[35]~combout ;
wire \cmd_mux_002|src_data[34]~combout ;
wire \cmd_mux_002|src_data[33]~combout ;
wire \cmd_mux_002|src_data[32]~combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_demux|src4_valid~0_combout ;
wire \cmd_demux|src4_valid~1_combout ;
wire \hps_h2f_lw_axi_master_rd_limiter|last_channel[4]~q ;
wire \cmd_demux_001|src4_valid~0_combout ;
wire \cmd_mux_004|src_valid~0_combout ;
wire \cmd_mux_004|src_valid~1_combout ;
wire \cmd_mux_004|src_payload[0]~combout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ;
wire \leds_s1_agent|cp_ready~0_combout ;
wire \leds_s1_agent|cp_ready~1_combout ;
wire \leds_s1_agent|uncompressor|last_packet_beat~2_combout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ;
wire \rsp_demux_004|WideOr0~0_combout ;
wire \leds_s1_agent_rsp_fifo|read~0_combout ;
wire \cmd_mux_004|src_data[78]~combout ;
wire \cmd_mux_004|src_data[79]~combout ;
wire \cmd_mux_004|src_data[35]~combout ;
wire \cmd_mux_004|src_data[34]~combout ;
wire \cmd_mux_004|src_data[33]~combout ;
wire \cmd_mux_004|src_data[32]~combout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ;
wire \cmd_demux|WideOr0~0_combout ;
wire \rsp_mux_001|src_payload~75_combout ;
wire \router|Equal3~8_combout ;
wire \control_s1_agent|rp_valid~combout ;
wire \base_address_ddr_s1_agent|rp_valid~combout ;
wire \leds_s1_agent|rp_valid~combout ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ;
wire \cmd_mux_003|src_payload~0_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector3~0_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector10~0_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector10~1_combout ;
wire \cmd_mux_003|src_data[73]~combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~0_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector4~1_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector11~1_combout ;
wire \cmd_mux_003|src_data[72]~combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~1_combout ;
wire \cmd_mux_003|src_payload~1_combout ;
wire \cmd_mux_003|src_payload~2_combout ;
wire \cmd_mux_003|src_payload~3_combout ;
wire \cmd_mux_003|src_payload~4_combout ;
wire \cmd_mux_003|src_payload~5_combout ;
wire \cmd_mux_003|src_payload~6_combout ;
wire \cmd_mux_003|src_payload~7_combout ;
wire \cmd_mux_003|src_payload~8_combout ;
wire \cmd_mux_003|src_payload~9_combout ;
wire \cmd_mux_003|src_payload~10_combout ;
wire \cmd_mux_003|src_payload~11_combout ;
wire \cmd_mux_003|src_payload~12_combout ;
wire \cmd_mux_003|src_payload~13_combout ;
wire \cmd_mux_003|src_payload~14_combout ;
wire \cmd_mux_003|src_payload~15_combout ;
wire \cmd_mux_003|src_payload~16_combout ;
wire \cmd_mux_003|src_payload~17_combout ;
wire \cmd_mux_003|src_payload~18_combout ;
wire \cmd_mux_003|src_payload~19_combout ;
wire \cmd_mux_003|src_payload~20_combout ;
wire \cmd_mux_003|src_payload~21_combout ;
wire \cmd_mux_003|src_payload~22_combout ;
wire \cmd_mux_003|src_payload~23_combout ;
wire \cmd_mux_003|src_payload~24_combout ;
wire \cmd_mux_003|src_payload~25_combout ;
wire \cmd_mux_003|src_payload~26_combout ;
wire \cmd_mux_003|src_payload~27_combout ;
wire \cmd_mux_003|src_payload~28_combout ;
wire \cmd_mux_003|src_payload~29_combout ;
wire \cmd_mux_003|src_payload~30_combout ;
wire \cmd_mux_003|src_payload~31_combout ;
wire \cmd_mux_002|src_payload~0_combout ;
wire \cmd_mux_002|src_data[73]~combout ;
wire \cmd_mux_002|src_data[72]~combout ;
wire \cmd_mux_002|src_payload~1_combout ;
wire \cmd_mux_002|src_payload~2_combout ;
wire \cmd_mux_002|src_payload~3_combout ;
wire \cmd_mux_002|src_payload~4_combout ;
wire \cmd_mux_002|src_payload~5_combout ;
wire \cmd_mux_002|src_payload~6_combout ;
wire \cmd_mux_002|src_payload~7_combout ;
wire \cmd_mux_002|src_payload~8_combout ;
wire \cmd_mux_002|src_payload~9_combout ;
wire \cmd_mux_002|src_payload~10_combout ;
wire \cmd_mux_002|src_payload~11_combout ;
wire \cmd_mux_002|src_payload~12_combout ;
wire \cmd_mux_002|src_payload~13_combout ;
wire \cmd_mux_002|src_payload~14_combout ;
wire \cmd_mux_002|src_payload~15_combout ;
wire \cmd_mux_002|src_payload~16_combout ;
wire \cmd_mux_002|src_payload~17_combout ;
wire \cmd_mux_002|src_payload~18_combout ;
wire \cmd_mux_002|src_payload~19_combout ;
wire \cmd_mux_002|src_payload~20_combout ;
wire \cmd_mux_002|src_payload~21_combout ;
wire \cmd_mux_002|src_payload~22_combout ;
wire \cmd_mux_002|src_payload~23_combout ;
wire \cmd_mux_002|src_payload~24_combout ;
wire \cmd_mux_002|src_payload~25_combout ;
wire \cmd_mux_002|src_payload~26_combout ;
wire \cmd_mux_002|src_payload~27_combout ;
wire \cmd_mux_002|src_payload~28_combout ;
wire \cmd_mux_002|src_payload~29_combout ;
wire \cmd_mux_002|src_payload~30_combout ;
wire \cmd_mux_002|src_payload~31_combout ;
wire \cmd_mux_004|src_payload~0_combout ;
wire \cmd_mux_004|src_data[73]~combout ;
wire \cmd_mux_004|src_data[72]~combout ;
wire \cmd_mux_004|src_payload~1_combout ;
wire \cmd_mux_004|src_payload~2_combout ;
wire \cmd_mux_004|src_payload~3_combout ;
wire \cmd_mux_004|src_payload~4_combout ;
wire \cmd_mux_004|src_payload~5_combout ;
wire \cmd_mux_004|src_payload~6_combout ;
wire \cmd_mux_004|src_payload~7_combout ;
wire \cmd_mux_004|src_payload~8_combout ;
wire \cmd_mux_004|src_payload~9_combout ;
wire \cmd_demux_001|WideOr0~1_combout ;
wire \router|Equal4~1_combout ;
wire \leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ;
wire \cmd_demux_001|src4_valid~1_combout ;
wire \cmd_mux_002|src_data[92]~combout ;
wire \cmd_mux_003|src_data[92]~combout ;
wire \cmd_mux_004|src_data[92]~combout ;
wire \cmd_mux_002|src_data[93]~combout ;
wire \cmd_mux_003|src_data[93]~combout ;
wire \cmd_mux_004|src_data[93]~combout ;
wire \cmd_mux_002|src_data[94]~combout ;
wire \cmd_mux_003|src_data[94]~combout ;
wire \cmd_mux_004|src_data[94]~combout ;
wire \cmd_mux_002|src_data[95]~combout ;
wire \cmd_mux_003|src_data[95]~combout ;
wire \cmd_mux_004|src_data[95]~combout ;
wire \cmd_mux_002|src_data[96]~combout ;
wire \cmd_mux_003|src_data[96]~combout ;
wire \cmd_mux_004|src_data[96]~combout ;
wire \cmd_mux_002|src_data[97]~combout ;
wire \cmd_mux_003|src_data[97]~combout ;
wire \cmd_mux_004|src_data[97]~combout ;
wire \cmd_mux_002|src_data[98]~combout ;
wire \cmd_mux_003|src_data[98]~combout ;
wire \cmd_mux_004|src_data[98]~combout ;
wire \cmd_mux_002|src_data[99]~combout ;
wire \cmd_mux_003|src_data[99]~combout ;
wire \cmd_mux_004|src_data[99]~combout ;
wire \cmd_mux_002|src_data[100]~combout ;
wire \cmd_mux_003|src_data[100]~combout ;
wire \cmd_mux_004|src_data[100]~combout ;
wire \cmd_mux_002|src_data[101]~combout ;
wire \cmd_mux_003|src_data[101]~combout ;
wire \cmd_mux_004|src_data[101]~combout ;
wire \cmd_mux_002|src_data[102]~combout ;
wire \cmd_mux_003|src_data[102]~combout ;
wire \cmd_mux_004|src_data[102]~combout ;
wire \cmd_mux_002|src_data[103]~combout ;
wire \cmd_mux_003|src_data[103]~combout ;
wire \cmd_mux_004|src_data[103]~combout ;
wire \cmd_mux_003|src_data[77]~combout ;
wire \cmd_mux_002|src_data[77]~combout ;
wire \cmd_mux_004|src_data[77]~combout ;
wire \cmd_mux|src_payload~0_combout ;
wire \cmd_mux|src_payload~1_combout ;
wire \cmd_mux|src_payload~2_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector5~1_combout ;
wire \hps_h2f_lw_axi_master_agent|Add3~3_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector12~0_combout ;
wire \cmd_mux_003|src_data[71]~combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~15_combout ;
wire \hps_h2f_lw_axi_master_agent|Decoder1~4_combout ;
wire \cmd_mux_002|src_data[71]~combout ;
wire \cmd_mux_004|src_data[71]~combout ;
wire \cmd_mux_001|src_payload~0_combout ;
wire \cmd_mux_001|src_payload~1_combout ;
wire \cmd_mux_001|src_payload~2_combout ;
wire \cmd_mux_005|src_payload~0_combout ;
wire \cmd_mux_005|src_payload~1_combout ;
wire \cmd_mux_005|src_payload~2_combout ;
wire \hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~16_combout ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ;
wire \hps_h2f_lw_axi_master_agent|Selector6~0_combout ;
wire \switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ;
wire \cmd_mux_003|src_data[70]~combout ;
wire \cmd_mux_002|src_data[70]~combout ;
wire \cmd_mux_004|src_data[70]~combout ;


terminal_qsys_altera_avalon_sc_fifo_6 rbf_id_control_slave_agent_rdata_fifo(
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.read_latency_shift_reg_0(\rbf_id_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\rbf_id_control_slave_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\rbf_id_control_slave_agent_rdata_fifo|empty~combout ),
	.mem_11_0(\rbf_id_control_slave_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_30(\rbf_id_control_slave_translator|av_readdata_pre[30]~q ),
	.mem_10_0(\rbf_id_control_slave_agent_rdata_fifo|mem[0][10]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.read(\rbf_id_control_slave_agent_rdata_fifo|read~0_combout ),
	.clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_7 rbf_id_control_slave_agent_rsp_fifo(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\rbf_id_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_60(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.wait_latency_counter_1(\rbf_id_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rbf_id_control_slave_translator|wait_latency_counter[0]~q ),
	.out_valid_reg(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_117_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][117]~q ),
	.mem_57_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_0(\rbf_id_control_slave_agent_rsp_fifo|mem_used[0]~q ),
	.mem_69_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][65]~q ),
	.mem_92_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][103]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.nxt_out_eop(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\rbf_id_control_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\rbf_id_control_slave_agent_rdata_fifo|read~0_combout ),
	.write(\rbf_id_control_slave_agent_rsp_fifo|write~0_combout ),
	.write1(\rbf_id_control_slave_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.in_data_reg_92(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_agent_3 rbf_id_control_slave_agent(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_data_reg_60(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_narrow_reg(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\rbf_id_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rbf_id_control_slave_translator|wait_latency_counter[0]~q ),
	.cp_ready(\rbf_id_control_slave_agent|cp_ready~0_combout ),
	.empty(\rbf_id_control_slave_agent_rdata_fifo|empty~combout ),
	.mem_57_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_0(\rbf_id_control_slave_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\rbf_id_control_slave_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\rbf_id_control_slave_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat1(\rbf_id_control_slave_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.last_packet_beat2(\rbf_id_control_slave_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\rbf_id_control_slave_agent_rdata_fifo|read~0_combout ),
	.cp_ready1(\rbf_id_control_slave_agent|cp_ready~1_combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_axi_master_ni hps_h2f_lw_axi_master_agent(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.h2f_lw_AWADDR_15(h2f_lw_AWADDR_15),
	.h2f_lw_AWADDR_16(h2f_lw_AWADDR_16),
	.h2f_lw_AWADDR_17(h2f_lw_AWADDR_17),
	.h2f_lw_AWADDR_18(h2f_lw_AWADDR_18),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_0(h2f_lw_AWLEN_0),
	.h2f_lw_AWLEN_1(h2f_lw_AWLEN_1),
	.h2f_lw_AWLEN_2(h2f_lw_AWLEN_2),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.address_burst_7(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_6(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.address_burst_9(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[9]~q ),
	.address_burst_8(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.address_burst_11(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[11]~q ),
	.address_burst_10(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[10]~q ),
	.address_burst_15(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[15]~q ),
	.address_burst_14(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[14]~q ),
	.address_burst_13(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[13]~q ),
	.address_burst_12(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[12]~q ),
	.Add5(\hps_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add51(\hps_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.write_addr_data_both_valid1(\hps_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ),
	.sop_enable1(\hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_5(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.address_burst_4(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[4]~q ),
	.out_data_18(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[18]~0_combout ),
	.out_data_17(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[17]~1_combout ),
	.out_data_16(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[16]~2_combout ),
	.nonposted_cmd_accepted(nonposted_cmd_accepted1),
	.Decoder1(\hps_h2f_lw_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out2),
	.burst_bytecount_6(\hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.burst_bytecount_5(\hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.burst_bytecount_4(\hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.burst_bytecount_3(\hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\hps_h2f_lw_axi_master_agent|write_cp_data[66]~3_combout ),
	.burst_bytecount_2(\hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\hps_h2f_lw_axi_master_agent|write_cp_data[65]~4_combout ),
	.Selector3(\hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_h2f_lw_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.base_address_3(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.Selector4(\hps_h2f_lw_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.base_address_2(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.Selector5(\hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Add3(\hps_h2f_lw_axi_master_agent|Add3~3_combout ),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.out_data_1(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~15_combout ),
	.Decoder11(\hps_h2f_lw_axi_master_agent|Decoder1~4_combout ),
	.out_data_0(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~16_combout ),
	.Selector6(\hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_slave_translator_5 switches_s1_translator(
	.wait_latency_counter_1(\switches_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\switches_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\switches_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\switches_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\switches_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\switches_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\switches_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\switches_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\switches_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\switches_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\switches_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\switches_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\switches_s1_translator|av_readdata_pre[9]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.write(\switches_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\switches_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_94,readdata_84,readdata_74,readdata_64,readdata_54,readdata_44,readdata_34,readdata_24,readdata_14,readdata_04}),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_translator_2 leds_s1_translator(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.out_valid_reg(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\leds_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.read_latency_shift_reg_0(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\leds_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\leds_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\leds_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\leds_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\leds_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\leds_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\leds_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\leds_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\leds_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\leds_s1_translator|av_readdata_pre[9]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.m0_write(m0_write2),
	.in_data_reg_60(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_93,readdata_82,readdata_72,readdata_62,readdata_52,readdata_42,readdata_32,readdata_22,readdata_12,readdata_02}),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_translator base_address_ddr_s1_translator(
	.out_valid_reg(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\base_address_ddr_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\base_address_ddr_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.read_latency_shift_reg_0(\base_address_ddr_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\base_address_ddr_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\base_address_ddr_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\base_address_ddr_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\base_address_ddr_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\base_address_ddr_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\base_address_ddr_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\base_address_ddr_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\base_address_ddr_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\base_address_ddr_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\base_address_ddr_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\base_address_ddr_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\base_address_ddr_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\base_address_ddr_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\base_address_ddr_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\base_address_ddr_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\base_address_ddr_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\base_address_ddr_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\base_address_ddr_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\base_address_ddr_s1_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\base_address_ddr_s1_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_20(\base_address_ddr_s1_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\base_address_ddr_s1_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\base_address_ddr_s1_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\base_address_ddr_s1_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\base_address_ddr_s1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\base_address_ddr_s1_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\base_address_ddr_s1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\base_address_ddr_s1_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\base_address_ddr_s1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\base_address_ddr_s1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\base_address_ddr_s1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\base_address_ddr_s1_translator|av_readdata_pre[31]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.m0_write(m0_write),
	.in_data_reg_60(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.av_readdata({readdata_311,readdata_301,readdata_29,readdata_281,readdata_271,readdata_26,readdata_25,readdata_242,readdata_231,readdata_221,readdata_212,readdata_201,readdata_191,readdata_18,readdata_17,readdata_16,readdata_15,readdata_141,readdata_131,readdata_121,readdata_112,
readdata_101,readdata_92,readdata_81,readdata_71,readdata_61,readdata_51,readdata_41,readdata_31,readdata_21,readdata_11,readdata_01}),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_translator_1 control_s1_translator(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.out_valid_reg(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\control_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\control_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.read_latency_shift_reg_0(\control_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\control_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\control_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\control_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\control_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\control_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\control_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\control_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\control_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\control_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\control_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\control_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\control_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\control_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\control_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\control_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\control_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\control_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\control_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\control_s1_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\control_s1_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_20(\control_s1_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\control_s1_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\control_s1_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\control_s1_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\control_s1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\control_s1_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\control_s1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\control_s1_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\control_s1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\control_s1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\control_s1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\control_s1_translator|av_readdata_pre[31]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.m0_write(m0_write1),
	.in_data_reg_60(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.av_readdata({readdata_312,readdata_30,readdata_291,readdata_28,readdata_27,readdata_261,readdata_251,readdata_241,readdata_232,readdata_222,readdata_211,readdata_20,readdata_19,readdata_181,readdata_171,readdata_161,readdata_151,readdata_142,readdata_132,readdata_122,readdata_111,
readdata_10,readdata_91,readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_translator_4 state_s1_translator(
	.wait_latency_counter_1(\state_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\state_s1_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\state_s1_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_0(\state_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_1(\state_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_2(\state_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_3(\state_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_4(\state_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_5(\state_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_6(\state_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\state_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_8(\state_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\state_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_10(\state_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_11(\state_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_12(\state_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_13(\state_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_14(\state_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\state_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_16(\state_s1_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_17(\state_s1_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_18(\state_s1_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_19(\state_s1_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_20(\state_s1_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_21(\state_s1_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_22(\state_s1_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_23(\state_s1_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_24(\state_s1_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_25(\state_s1_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_26(\state_s1_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_27(\state_s1_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_28(\state_s1_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_29(\state_s1_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_30(\state_s1_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_31(\state_s1_translator|av_readdata_pre[31]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(\state_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\state_s1_agent_rsp_fifo|write~1_combout ),
	.av_readdata({readdata_313,readdata_302,readdata_292,readdata_282,readdata_272,readdata_262,readdata_252,readdata_243,readdata_233,readdata_223,readdata_213,readdata_202,readdata_192,readdata_182,readdata_172,readdata_162,readdata_152,readdata_143,readdata_133,readdata_123,readdata_113,
readdata_102,readdata_9,readdata_83,readdata_73,readdata_63,readdata_53,readdata_43,readdata_33,readdata_23,readdata_13,readdata_03}),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_translator_3 rbf_id_control_slave_translator(
	.wait_latency_counter_1(\rbf_id_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\rbf_id_control_slave_translator|wait_latency_counter[0]~q ),
	.read_latency_shift_reg_0(\rbf_id_control_slave_translator|read_latency_shift_reg[0]~q ),
	.av_readdata_pre_30(\rbf_id_control_slave_translator|av_readdata_pre[30]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.write(\rbf_id_control_slave_agent_rsp_fifo|write~0_combout ),
	.write1(\rbf_id_control_slave_agent_rsp_fifo|write~1_combout ),
	.av_readdata({gnd,\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.clk(clk_clk));

terminal_qsys_altera_merlin_burst_adapter_1 control_s1_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.nxt_in_ready(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_narrow_reg(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_59(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.write(\control_s1_agent_rsp_fifo|write~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.sop_enable(\hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal31(\router|Equal3~7_combout ),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.in_data_reg_0(in_data_reg_01),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_31),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_21),
	.in_data_reg_1(in_data_reg_110),
	.in_data_reg_2(in_data_reg_210),
	.in_data_reg_3(in_data_reg_32),
	.in_data_reg_4(in_data_reg_41),
	.in_data_reg_5(in_data_reg_51),
	.in_data_reg_6(in_data_reg_61),
	.in_data_reg_7(in_data_reg_71),
	.in_data_reg_8(in_data_reg_81),
	.in_data_reg_9(in_data_reg_91),
	.in_data_reg_10(in_data_reg_101),
	.in_data_reg_11(in_data_reg_111),
	.in_data_reg_12(in_data_reg_121),
	.in_data_reg_13(in_data_reg_131),
	.in_data_reg_14(in_data_reg_141),
	.in_data_reg_15(in_data_reg_151),
	.in_data_reg_16(in_data_reg_161),
	.in_data_reg_17(in_data_reg_171),
	.in_data_reg_18(in_data_reg_181),
	.in_data_reg_19(in_data_reg_191),
	.in_data_reg_20(in_data_reg_201),
	.in_data_reg_21(in_data_reg_211),
	.in_data_reg_22(in_data_reg_221),
	.in_data_reg_23(in_data_reg_231),
	.in_data_reg_24(in_data_reg_241),
	.in_data_reg_25(in_data_reg_251),
	.in_data_reg_26(in_data_reg_261),
	.in_data_reg_27(in_data_reg_271),
	.in_data_reg_28(in_data_reg_281),
	.in_data_reg_29(in_data_reg_291),
	.in_data_reg_30(in_data_reg_301),
	.in_data_reg_31(in_data_reg_311),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.burst_bytecount_6(\hps_h2f_lw_axi_master_agent|burst_bytecount[6]~q ),
	.write_cp_data_69(\hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.burst_bytecount_5(\hps_h2f_lw_axi_master_agent|burst_bytecount[5]~q ),
	.write_cp_data_68(\hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.burst_bytecount_4(\hps_h2f_lw_axi_master_agent|burst_bytecount[4]~q ),
	.write_cp_data_67(\hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.burst_bytecount_3(\hps_h2f_lw_axi_master_agent|burst_bytecount[3]~q ),
	.write_cp_data_66(\hps_h2f_lw_axi_master_agent|write_cp_data[66]~3_combout ),
	.burst_bytecount_2(\hps_h2f_lw_axi_master_agent|burst_bytecount[2]~q ),
	.write_cp_data_65(\hps_h2f_lw_axi_master_agent|write_cp_data[65]~4_combout ),
	.WideNor0(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src_valid(\cmd_mux_002|src_valid~0_combout ),
	.src_payload_0(\cmd_mux_002|src_payload[0]~combout ),
	.nxt_out_eop(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready(\control_s1_agent|cp_ready~2_combout ),
	.in_data_reg_60(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux_002|src_data[78]~combout ),
	.src_data_79(\cmd_mux_002|src_data[79]~combout ),
	.src_data_35(\cmd_mux_002|src_data[35]~combout ),
	.src_data_34(\cmd_mux_002|src_data[34]~combout ),
	.src_data_33(\cmd_mux_002|src_data[33]~combout ),
	.src_data_32(\cmd_mux_002|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_6(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_92(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.base_address_3(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.base_address_2(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_002|src_payload~0_combout ),
	.src_data_73(\cmd_mux_002|src_data[73]~combout ),
	.src_data_72(\cmd_mux_002|src_data[72]~combout ),
	.src_payload1(\cmd_mux_002|src_payload~1_combout ),
	.src_payload2(\cmd_mux_002|src_payload~2_combout ),
	.src_payload3(\cmd_mux_002|src_payload~3_combout ),
	.src_payload4(\cmd_mux_002|src_payload~4_combout ),
	.src_payload5(\cmd_mux_002|src_payload~5_combout ),
	.src_payload6(\cmd_mux_002|src_payload~6_combout ),
	.src_payload7(\cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\cmd_mux_002|src_payload~31_combout ),
	.src_data_92(\cmd_mux_002|src_data[92]~combout ),
	.src_data_93(\cmd_mux_002|src_data[93]~combout ),
	.src_data_94(\cmd_mux_002|src_data[94]~combout ),
	.src_data_95(\cmd_mux_002|src_data[95]~combout ),
	.src_data_96(\cmd_mux_002|src_data[96]~combout ),
	.src_data_97(\cmd_mux_002|src_data[97]~combout ),
	.src_data_98(\cmd_mux_002|src_data[98]~combout ),
	.src_data_99(\cmd_mux_002|src_data[99]~combout ),
	.src_data_100(\cmd_mux_002|src_data[100]~combout ),
	.src_data_101(\cmd_mux_002|src_data[101]~combout ),
	.src_data_102(\cmd_mux_002|src_data[102]~combout ),
	.src_data_103(\cmd_mux_002|src_data[103]~combout ),
	.src_data_77(\cmd_mux_002|src_data[77]~combout ),
	.out_data_1(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~15_combout ),
	.src_data_71(\cmd_mux_002|src_data[71]~combout ),
	.out_data_0(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~16_combout ),
	.src_data_70(\cmd_mux_002|src_data[70]~combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_burst_adapter_4 state_s1_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\state_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_60(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_narrow_reg(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\state_s1_agent|cp_ready~0_combout ),
	.nxt_in_ready(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(\hps_h2f_lw_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.nxt_out_eop(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.Equal2(\router_001|Equal2~0_combout ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.src_valid1(\cmd_mux_001|src_valid~1_combout ),
	.out_byte_cnt_reg_2(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready1(\state_s1_agent|cp_ready~1_combout ),
	.out_uncomp_byte_cnt_reg_5(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_92(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.Selector10(\hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_33),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_23),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_payload1(\cmd_mux_001|src_payload~1_combout ),
	.src_payload2(\cmd_mux_001|src_payload~2_combout ),
	.nxt_out_burstwrap_1(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_out_burstwrap_0(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_burst_adapter_3 rbf_id_control_slave_burst_adapter(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.has_pending_responses(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.stateST_COMP_TRANS(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\rbf_id_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_60(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_narrow_reg(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\rbf_id_control_slave_agent|cp_ready~0_combout ),
	.nxt_in_ready(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.Decoder1(\hps_h2f_lw_axi_master_agent|Decoder1~0_combout ),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.nxt_out_eop(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.Equal1(\router_001|Equal1~3_combout ),
	.last_channel_0(\hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.out_byte_cnt_reg_2(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.cp_ready1(\rbf_id_control_slave_agent|cp_ready~1_combout ),
	.out_uncomp_byte_cnt_reg_6(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.out_uncomp_byte_cnt_reg_5(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.int_nxt_addr_reg_dly_2(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|int_nxt_addr_reg_dly[2]~q ),
	.in_data_reg_92(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.nxt_out_burstwrap_1(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_out_burstwrap_0(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_traffic_limiter hps_h2f_lw_axi_master_rd_limiter(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.h2f_lw_ARADDR_16(h2f_lw_ARADDR_16),
	.h2f_lw_ARADDR_17(h2f_lw_ARADDR_17),
	.h2f_lw_ARADDR_18(h2f_lw_ARADDR_18),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.cmd_sink_channel({\router_001|Equal5~0_combout ,\router_001|src_channel[4]~1_combout ,\router_001|Equal4~1_combout ,\router_001|Equal3~0_combout ,\router_001|Equal2~0_combout ,\router_001|Equal1~3_combout }),
	.sink_ready(\cmd_demux_001|sink_ready~0_combout ),
	.has_pending_responses1(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router_001|src_data[91]~1_combout ,\router_001|src_data[90]~0_combout ,\router_001|src_channel[4]~0_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.sink_ready1(\cmd_demux_001|sink_ready~1_combout ),
	.WideOr0(\cmd_demux_001|WideOr0~0_combout ),
	.sink_ready2(\cmd_demux_001|sink_ready~4_combout ),
	.sink_ready3(\cmd_demux_001|sink_ready~5_combout ),
	.cmd_sink_ready(cmd_sink_ready),
	.src_payload_0(src_payload_0),
	.WideOr1(WideOr11),
	.last_channel_5(\hps_h2f_lw_axi_master_rd_limiter|last_channel[5]~q ),
	.WideOr01(\cmd_demux_001|WideOr0~combout ),
	.reset(altera_reset_synchronizer_int_chain_out2),
	.last_channel_3(\hps_h2f_lw_axi_master_rd_limiter|last_channel[3]~q ),
	.last_channel_0(\hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ),
	.last_channel_1(\hps_h2f_lw_axi_master_rd_limiter|last_channel[1]~q ),
	.last_channel_2(\hps_h2f_lw_axi_master_rd_limiter|last_channel[2]~q ),
	.last_channel_4(\hps_h2f_lw_axi_master_rd_limiter|last_channel[4]~q ),
	.WideOr02(\cmd_demux_001|WideOr0~1_combout ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_traffic_limiter_1 hps_h2f_lw_axi_master_wr_limiter(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.write_addr_data_both_valid(\hps_h2f_lw_axi_master_agent|write_addr_data_both_valid~combout ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal31(\router|Equal3~7_combout ),
	.Equal4(\router|Equal4~0_combout ),
	.has_pending_responses1(\hps_h2f_lw_axi_master_wr_limiter|has_pending_responses~q ),
	.last_channel_2(\hps_h2f_lw_axi_master_wr_limiter|last_channel[2]~q ),
	.last_channel_4(\hps_h2f_lw_axi_master_wr_limiter|last_channel[4]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ),
	.sink_ready2(\cmd_demux|sink_ready~2_combout ),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.src0_valid(\rsp_demux_002|src0_valid~combout ),
	.mem_57_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux_003|src0_valid~combout ),
	.mem_57_01(\leds_s1_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid2(\rsp_demux_004|src0_valid~combout ),
	.WideOr1(WideOr1),
	.comb(\base_address_ddr_s1_agent|comb~0_combout ),
	.mem_117_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][117]~q ),
	.last_packet_beat(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb1(\leds_s1_agent|comb~0_combout ),
	.mem_117_01(\leds_s1_agent_rsp_fifo|mem[0][117]~q ),
	.last_packet_beat2(\leds_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat3(\leds_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted1),
	.reset(altera_reset_synchronizer_int_chain_out2),
	.last_channel_3(\hps_h2f_lw_axi_master_wr_limiter|last_channel[3]~q ),
	.cmd_sink_channel({gnd,\cmd_demux|src4_valid~0_combout ,\router|Equal4~1_combout ,\router|Equal3~8_combout ,gnd,gnd}),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.src_payload(\rsp_mux_001|src_payload~75_combout ),
	.clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_router_1 router_001(
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_4(h2f_lw_ARADDR_4),
	.h2f_lw_ARADDR_5(h2f_lw_ARADDR_5),
	.h2f_lw_ARADDR_6(h2f_lw_ARADDR_6),
	.h2f_lw_ARADDR_7(h2f_lw_ARADDR_7),
	.h2f_lw_ARADDR_8(h2f_lw_ARADDR_8),
	.h2f_lw_ARADDR_9(h2f_lw_ARADDR_9),
	.h2f_lw_ARADDR_10(h2f_lw_ARADDR_10),
	.h2f_lw_ARADDR_11(h2f_lw_ARADDR_11),
	.h2f_lw_ARADDR_12(h2f_lw_ARADDR_12),
	.h2f_lw_ARADDR_13(h2f_lw_ARADDR_13),
	.h2f_lw_ARADDR_14(h2f_lw_ARADDR_14),
	.h2f_lw_ARADDR_15(h2f_lw_ARADDR_15),
	.h2f_lw_ARADDR_16(h2f_lw_ARADDR_16),
	.h2f_lw_ARADDR_17(h2f_lw_ARADDR_17),
	.h2f_lw_ARADDR_18(h2f_lw_ARADDR_18),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.Equal5(\router_001|Equal5~0_combout ),
	.src_channel_4(\router_001|src_channel[4]~0_combout ),
	.Equal4(\router_001|Equal4~0_combout ),
	.Equal41(\router_001|Equal4~1_combout ),
	.Equal12(\router_001|Equal1~2_combout ),
	.Equal3(\router_001|Equal3~0_combout ),
	.src_channel_41(\router_001|src_channel[4]~1_combout ),
	.src_data_90(\router_001|src_data[90]~0_combout ),
	.src_data_91(\router_001|src_data[91]~1_combout ),
	.Equal13(\router_001|Equal1~3_combout ),
	.Equal2(\router_001|Equal2~0_combout ));

terminal_qsys_terminal_qsys_mm_interconnect_0_router router(
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.h2f_lw_AWADDR_15(h2f_lw_AWADDR_15),
	.address_burst_7(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[7]~q ),
	.address_burst_6(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[6]~q ),
	.address_burst_9(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[9]~q ),
	.address_burst_8(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[8]~q ),
	.address_burst_11(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[11]~q ),
	.address_burst_10(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[10]~q ),
	.address_burst_15(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[15]~q ),
	.address_burst_14(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[14]~q ),
	.address_burst_13(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[13]~q ),
	.address_burst_12(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[12]~q ),
	.sop_enable(\hps_h2f_lw_axi_master_agent|sop_enable~q ),
	.address_burst_5(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[5]~q ),
	.address_burst_4(\hps_h2f_lw_axi_master_agent|align_address_to_size|address_burst[4]~q ),
	.Equal3(\router|Equal3~6_combout ),
	.out_data_18(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[18]~0_combout ),
	.out_data_17(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[17]~1_combout ),
	.out_data_16(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[16]~2_combout ),
	.Equal31(\router|Equal3~7_combout ),
	.Equal4(\router|Equal4~0_combout ),
	.Equal32(\router|Equal3~8_combout ),
	.Equal41(\router|Equal4~1_combout ));

terminal_qsys_altera_avalon_sc_fifo_10 switches_s1_agent_rdata_fifo(
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\switches_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\switches_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\switches_s1_agent_rdata_fifo|empty~combout ),
	.mem_0_0(\switches_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_0(\switches_s1_translator|av_readdata_pre[0]~q ),
	.mem_1_0(\switches_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_1(\switches_s1_translator|av_readdata_pre[1]~q ),
	.mem_2_0(\switches_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_2(\switches_s1_translator|av_readdata_pre[2]~q ),
	.mem_3_0(\switches_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_3(\switches_s1_translator|av_readdata_pre[3]~q ),
	.mem_4_0(\switches_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_4(\switches_s1_translator|av_readdata_pre[4]~q ),
	.mem_5_0(\switches_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_5(\switches_s1_translator|av_readdata_pre[5]~q ),
	.mem_6_0(\switches_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_6(\switches_s1_translator|av_readdata_pre[6]~q ),
	.mem_7_0(\switches_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_7(\switches_s1_translator|av_readdata_pre[7]~q ),
	.mem_8_0(\switches_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_8(\switches_s1_translator|av_readdata_pre[8]~q ),
	.mem_9_0(\switches_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_9(\switches_s1_translator|av_readdata_pre[9]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.read(\switches_s1_agent_rdata_fifo|read~0_combout ),
	.clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_11 switches_s1_agent_rsp_fifo(
	.mem_used_1(\switches_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_60(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.wait_latency_counter_1(\switches_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\switches_s1_translator|wait_latency_counter[0]~q ),
	.out_valid_reg(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_117_0(\switches_s1_agent_rsp_fifo|mem[0][117]~q ),
	.mem_57_0(\switches_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_0(\switches_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_69_0(\switches_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\switches_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\switches_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\switches_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\switches_s1_agent_rsp_fifo|mem[0][65]~q ),
	.mem_92_0(\switches_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\switches_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\switches_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\switches_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\switches_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\switches_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\switches_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\switches_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\switches_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\switches_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\switches_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\switches_s1_agent_rsp_fifo|mem[0][103]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.nxt_out_eop(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\switches_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\switches_s1_agent_rdata_fifo|read~0_combout ),
	.write(\switches_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\switches_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_92(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_agent_5 switches_s1_agent(
	.stateST_COMP_TRANS(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_data_reg_60(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_narrow_reg(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\switches_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\switches_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\switches_s1_agent|cp_ready~0_combout ),
	.empty(\switches_s1_agent_rdata_fifo|empty~combout ),
	.mem_57_0(\switches_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_0(\switches_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\switches_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\switches_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\switches_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\switches_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\switches_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\switches_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat1(\switches_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.last_packet_beat2(\switches_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\switches_s1_agent_rdata_fifo|read~0_combout ),
	.cp_ready1(\switches_s1_agent|cp_ready~1_combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_4 leds_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\leds_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\leds_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\leds_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\leds_s1_translator|av_readdata_pre[0]~q ),
	.always4(\leds_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\leds_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\leds_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\leds_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\leds_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\leds_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\leds_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\leds_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\leds_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\leds_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\leds_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\leds_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\leds_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\leds_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\leds_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\leds_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_8(\leds_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\leds_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_9(\leds_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\leds_s1_agent_rdata_fifo|mem[0][9]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.WideOr0(\rsp_demux_004|WideOr0~0_combout ),
	.clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_5 leds_s1_agent_rsp_fifo(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.out_valid_reg(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\leds_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.in_data_reg_59(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.local_write(\leds_s1_agent|local_write~combout ),
	.write(\leds_s1_agent_rsp_fifo|write~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_116_0(\leds_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_0(\leds_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\leds_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\leds_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\leds_s1_agent|comb~0_combout ),
	.mem_117_0(\leds_s1_agent_rsp_fifo|mem[0][117]~q ),
	.mem_69_0(\leds_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\leds_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\leds_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\leds_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\leds_s1_agent_rsp_fifo|mem[0][65]~q ),
	.mem_92_0(\leds_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\leds_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\leds_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\leds_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\leds_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\leds_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\leds_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\leds_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\leds_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\leds_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\leds_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\leds_s1_agent_rsp_fifo|mem[0][103]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.nxt_out_eop(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\leds_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.in_data_reg_60(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.WideOr01(\rsp_demux_004|WideOr0~0_combout ),
	.read(\leds_s1_agent_rsp_fifo|read~0_combout ),
	.out_byte_cnt_reg_2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_3(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_6(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.rp_valid(\leds_s1_agent|rp_valid~combout ),
	.in_data_reg_92(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_agent_2 leds_s1_agent(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\leds_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_12),
	.wait_latency_counter_0(wait_latency_counter_02),
	.in_data_reg_59(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.local_write1(\leds_s1_agent|local_write~combout ),
	.read_latency_shift_reg_0(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\leds_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\leds_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\leds_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_57_0(\leds_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\leds_s1_agent|comb~0_combout ),
	.last_packet_beat(\leds_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\leds_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\leds_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\leds_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\leds_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\leds_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat1(\leds_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.m0_write1(m0_write2),
	.cp_ready(\leds_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\leds_s1_agent|cp_ready~1_combout ),
	.last_packet_beat2(\leds_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\leds_s1_agent_rsp_fifo|read~0_combout ),
	.rp_valid1(\leds_s1_agent|rp_valid~combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo base_address_ddr_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\base_address_ddr_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\base_address_ddr_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\base_address_ddr_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\base_address_ddr_s1_translator|av_readdata_pre[0]~q ),
	.always4(\base_address_ddr_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\base_address_ddr_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\base_address_ddr_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\base_address_ddr_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\base_address_ddr_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\base_address_ddr_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\base_address_ddr_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\base_address_ddr_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_8(\base_address_ddr_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_9(\base_address_ddr_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_10(\base_address_ddr_s1_translator|av_readdata_pre[10]~q ),
	.mem_10_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_11(\base_address_ddr_s1_translator|av_readdata_pre[11]~q ),
	.mem_11_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_12(\base_address_ddr_s1_translator|av_readdata_pre[12]~q ),
	.mem_12_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_13(\base_address_ddr_s1_translator|av_readdata_pre[13]~q ),
	.mem_13_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_14(\base_address_ddr_s1_translator|av_readdata_pre[14]~q ),
	.mem_14_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_15(\base_address_ddr_s1_translator|av_readdata_pre[15]~q ),
	.mem_15_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_16(\base_address_ddr_s1_translator|av_readdata_pre[16]~q ),
	.mem_16_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_17(\base_address_ddr_s1_translator|av_readdata_pre[17]~q ),
	.mem_17_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_18(\base_address_ddr_s1_translator|av_readdata_pre[18]~q ),
	.mem_18_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_19(\base_address_ddr_s1_translator|av_readdata_pre[19]~q ),
	.mem_19_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_20(\base_address_ddr_s1_translator|av_readdata_pre[20]~q ),
	.mem_20_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_21(\base_address_ddr_s1_translator|av_readdata_pre[21]~q ),
	.mem_21_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_22(\base_address_ddr_s1_translator|av_readdata_pre[22]~q ),
	.mem_22_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_23(\base_address_ddr_s1_translator|av_readdata_pre[23]~q ),
	.mem_23_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_24(\base_address_ddr_s1_translator|av_readdata_pre[24]~q ),
	.mem_24_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_25(\base_address_ddr_s1_translator|av_readdata_pre[25]~q ),
	.mem_25_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_26(\base_address_ddr_s1_translator|av_readdata_pre[26]~q ),
	.mem_26_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_27(\base_address_ddr_s1_translator|av_readdata_pre[27]~q ),
	.mem_27_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_28(\base_address_ddr_s1_translator|av_readdata_pre[28]~q ),
	.mem_28_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_29(\base_address_ddr_s1_translator|av_readdata_pre[29]~q ),
	.mem_29_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_30(\base_address_ddr_s1_translator|av_readdata_pre[30]~q ),
	.mem_30_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_31(\base_address_ddr_s1_translator|av_readdata_pre[31]~q ),
	.mem_31_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][31]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.WideOr0(\rsp_demux_003|WideOr0~0_combout ),
	.clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_1 base_address_ddr_s1_agent_rsp_fifo(
	.out_valid_reg(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\base_address_ddr_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\base_address_ddr_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_59(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.local_write(\base_address_ddr_s1_agent|local_write~combout ),
	.write(\base_address_ddr_s1_agent_rsp_fifo|write~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_116_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_0(\base_address_ddr_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\base_address_ddr_s1_agent|comb~0_combout ),
	.mem_117_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][117]~q ),
	.mem_69_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][65]~q ),
	.mem_92_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][103]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.in_data_reg_60(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.WideOr01(\rsp_demux_003|WideOr0~0_combout ),
	.read(\base_address_ddr_s1_agent_rsp_fifo|read~0_combout ),
	.out_byte_cnt_reg_2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.rp_valid(\base_address_ddr_s1_agent|rp_valid~combout ),
	.in_data_reg_92(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_agent base_address_ddr_s1_agent(
	.stateST_COMP_TRANS(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\base_address_ddr_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\base_address_ddr_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.in_data_reg_59(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.local_write1(\base_address_ddr_s1_agent|local_write~combout ),
	.read_latency_shift_reg_0(\base_address_ddr_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\base_address_ddr_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\base_address_ddr_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_57_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\base_address_ddr_s1_agent|comb~0_combout ),
	.last_packet_beat(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat1(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.m0_write1(m0_write),
	.cp_ready(\base_address_ddr_s1_agent|cp_ready~2_combout ),
	.last_packet_beat2(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\base_address_ddr_s1_agent_rsp_fifo|read~0_combout ),
	.rp_valid1(\base_address_ddr_s1_agent|rp_valid~combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_2 control_s1_agent_rdata_fifo(
	.read_latency_shift_reg_0(\control_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\control_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\control_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\control_s1_agent_rsp_fifo|mem_used[0]~q ),
	.av_readdata_pre_0(\control_s1_translator|av_readdata_pre[0]~q ),
	.always4(\control_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\control_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_1(\control_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\control_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_2(\control_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\control_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_3(\control_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\control_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_4(\control_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\control_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_5(\control_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\control_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_6(\control_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\control_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_7(\control_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\control_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_8(\control_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\control_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_9(\control_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\control_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_10(\control_s1_translator|av_readdata_pre[10]~q ),
	.mem_10_0(\control_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_11(\control_s1_translator|av_readdata_pre[11]~q ),
	.mem_11_0(\control_s1_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_12(\control_s1_translator|av_readdata_pre[12]~q ),
	.mem_12_0(\control_s1_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_13(\control_s1_translator|av_readdata_pre[13]~q ),
	.mem_13_0(\control_s1_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_14(\control_s1_translator|av_readdata_pre[14]~q ),
	.mem_14_0(\control_s1_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_15(\control_s1_translator|av_readdata_pre[15]~q ),
	.mem_15_0(\control_s1_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_16(\control_s1_translator|av_readdata_pre[16]~q ),
	.mem_16_0(\control_s1_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_17(\control_s1_translator|av_readdata_pre[17]~q ),
	.mem_17_0(\control_s1_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_18(\control_s1_translator|av_readdata_pre[18]~q ),
	.mem_18_0(\control_s1_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_19(\control_s1_translator|av_readdata_pre[19]~q ),
	.mem_19_0(\control_s1_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_20(\control_s1_translator|av_readdata_pre[20]~q ),
	.mem_20_0(\control_s1_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_21(\control_s1_translator|av_readdata_pre[21]~q ),
	.mem_21_0(\control_s1_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_22(\control_s1_translator|av_readdata_pre[22]~q ),
	.mem_22_0(\control_s1_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_23(\control_s1_translator|av_readdata_pre[23]~q ),
	.mem_23_0(\control_s1_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_24(\control_s1_translator|av_readdata_pre[24]~q ),
	.mem_24_0(\control_s1_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_25(\control_s1_translator|av_readdata_pre[25]~q ),
	.mem_25_0(\control_s1_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_26(\control_s1_translator|av_readdata_pre[26]~q ),
	.mem_26_0(\control_s1_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_27(\control_s1_translator|av_readdata_pre[27]~q ),
	.mem_27_0(\control_s1_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_28(\control_s1_translator|av_readdata_pre[28]~q ),
	.mem_28_0(\control_s1_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_29(\control_s1_translator|av_readdata_pre[29]~q ),
	.mem_29_0(\control_s1_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_30(\control_s1_translator|av_readdata_pre[30]~q ),
	.mem_30_0(\control_s1_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_31(\control_s1_translator|av_readdata_pre[31]~q ),
	.mem_31_0(\control_s1_agent_rdata_fifo|mem[0][31]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.WideOr0(\rsp_demux_002|WideOr0~0_combout ),
	.clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_3 control_s1_agent_rsp_fifo(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.out_valid_reg(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\control_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\control_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.in_data_reg_59(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.local_write(\control_s1_agent|local_write~combout ),
	.write(\control_s1_agent_rsp_fifo|write~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_116_0(\control_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_0(\control_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\control_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\control_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\control_s1_agent|comb~0_combout ),
	.mem_117_0(\control_s1_agent_rsp_fifo|mem[0][117]~q ),
	.mem_69_0(\control_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\control_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\control_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\control_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\control_s1_agent_rsp_fifo|mem[0][65]~q ),
	.mem_92_0(\control_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\control_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\control_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\control_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\control_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\control_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\control_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\control_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\control_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\control_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\control_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\control_s1_agent_rsp_fifo|mem[0][103]~q ),
	.reset(altera_reset_synchronizer_int_chain_out1),
	.nxt_out_eop(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\control_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.in_data_reg_60(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.WideOr01(\rsp_demux_002|WideOr0~0_combout ),
	.read(\control_s1_agent_rsp_fifo|read~0_combout ),
	.out_byte_cnt_reg_2(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_3(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_6(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.rp_valid(\control_s1_agent|rp_valid~combout ),
	.in_data_reg_92(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_agent_1 control_s1_agent(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\control_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.WideOr0(\control_s1_agent|WideOr0~0_combout ),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.in_data_reg_59(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.local_write1(\control_s1_agent|local_write~combout ),
	.read_latency_shift_reg_0(\control_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\control_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\control_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\control_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_57_0(\control_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\control_s1_agent|comb~0_combout ),
	.last_packet_beat(\control_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\control_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\control_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\control_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\control_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\control_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat1(\control_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.m0_write1(m0_write1),
	.cp_ready(\control_s1_agent|cp_ready~2_combout ),
	.last_packet_beat2(\control_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\control_s1_agent_rsp_fifo|read~0_combout ),
	.rp_valid1(\control_s1_agent|rp_valid~combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_8 state_s1_agent_rdata_fifo(
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\state_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\state_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\state_s1_agent_rdata_fifo|empty~combout ),
	.mem_0_0(\state_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_0(\state_s1_translator|av_readdata_pre[0]~q ),
	.mem_1_0(\state_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_1(\state_s1_translator|av_readdata_pre[1]~q ),
	.mem_2_0(\state_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_2(\state_s1_translator|av_readdata_pre[2]~q ),
	.mem_3_0(\state_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_3(\state_s1_translator|av_readdata_pre[3]~q ),
	.mem_4_0(\state_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_4(\state_s1_translator|av_readdata_pre[4]~q ),
	.mem_5_0(\state_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_5(\state_s1_translator|av_readdata_pre[5]~q ),
	.mem_6_0(\state_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_6(\state_s1_translator|av_readdata_pre[6]~q ),
	.mem_7_0(\state_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_7(\state_s1_translator|av_readdata_pre[7]~q ),
	.mem_8_0(\state_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_8(\state_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_9(\state_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\state_s1_agent_rdata_fifo|mem[0][9]~q ),
	.mem_10_0(\state_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_10(\state_s1_translator|av_readdata_pre[10]~q ),
	.mem_11_0(\state_s1_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_11(\state_s1_translator|av_readdata_pre[11]~q ),
	.mem_12_0(\state_s1_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_12(\state_s1_translator|av_readdata_pre[12]~q ),
	.mem_13_0(\state_s1_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_13(\state_s1_translator|av_readdata_pre[13]~q ),
	.mem_14_0(\state_s1_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_14(\state_s1_translator|av_readdata_pre[14]~q ),
	.mem_15_0(\state_s1_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_15(\state_s1_translator|av_readdata_pre[15]~q ),
	.mem_16_0(\state_s1_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_16(\state_s1_translator|av_readdata_pre[16]~q ),
	.mem_17_0(\state_s1_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_17(\state_s1_translator|av_readdata_pre[17]~q ),
	.mem_18_0(\state_s1_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_18(\state_s1_translator|av_readdata_pre[18]~q ),
	.mem_19_0(\state_s1_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_19(\state_s1_translator|av_readdata_pre[19]~q ),
	.mem_20_0(\state_s1_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_20(\state_s1_translator|av_readdata_pre[20]~q ),
	.mem_21_0(\state_s1_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_21(\state_s1_translator|av_readdata_pre[21]~q ),
	.mem_22_0(\state_s1_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_22(\state_s1_translator|av_readdata_pre[22]~q ),
	.mem_23_0(\state_s1_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_23(\state_s1_translator|av_readdata_pre[23]~q ),
	.mem_24_0(\state_s1_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_24(\state_s1_translator|av_readdata_pre[24]~q ),
	.mem_25_0(\state_s1_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_25(\state_s1_translator|av_readdata_pre[25]~q ),
	.mem_26_0(\state_s1_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_26(\state_s1_translator|av_readdata_pre[26]~q ),
	.mem_27_0(\state_s1_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_27(\state_s1_translator|av_readdata_pre[27]~q ),
	.mem_28_0(\state_s1_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_28(\state_s1_translator|av_readdata_pre[28]~q ),
	.mem_29_0(\state_s1_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_29(\state_s1_translator|av_readdata_pre[29]~q ),
	.mem_30_0(\state_s1_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_30(\state_s1_translator|av_readdata_pre[30]~q ),
	.mem_31_0(\state_s1_agent_rdata_fifo|mem[0][31]~q ),
	.av_readdata_pre_31(\state_s1_translator|av_readdata_pre[31]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read(\state_s1_agent_rdata_fifo|read~0_combout ),
	.clk(clk_clk));

terminal_qsys_altera_avalon_sc_fifo_9 state_s1_agent_rsp_fifo(
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_used_1(\state_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_60(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.wait_latency_counter_1(\state_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\state_s1_translator|wait_latency_counter[0]~q ),
	.out_valid_reg(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.mem_117_0(\state_s1_agent_rsp_fifo|mem[0][117]~q ),
	.mem_57_0(\state_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_0(\state_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_69_0(\state_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\state_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\state_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\state_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\state_s1_agent_rsp_fifo|mem[0][65]~q ),
	.mem_92_0(\state_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\state_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\state_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\state_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\state_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\state_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\state_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\state_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\state_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\state_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\state_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\state_s1_agent_rsp_fifo|mem[0][103]~q ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_packet_beat(\state_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\state_s1_agent_rdata_fifo|read~0_combout ),
	.write(\state_s1_agent_rsp_fifo|write~0_combout ),
	.write1(\state_s1_agent_rsp_fifo|write~1_combout ),
	.out_byte_cnt_reg_2(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_92(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.clk(clk_clk));

terminal_qsys_altera_merlin_slave_agent_4 state_s1_agent(
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.stateST_COMP_TRANS(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.in_data_reg_60(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_narrow_reg(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.wait_latency_counter_1(\state_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\state_s1_translator|wait_latency_counter[0]~q ),
	.cp_ready(\state_s1_agent|cp_ready~0_combout ),
	.empty(\state_s1_agent_rdata_fifo|empty~combout ),
	.mem_57_0(\state_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_0(\state_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat(\state_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.mem_69_0(\state_s1_agent_rsp_fifo|mem[0][69]~q ),
	.mem_68_0(\state_s1_agent_rsp_fifo|mem[0][68]~q ),
	.mem_67_0(\state_s1_agent_rsp_fifo|mem[0][67]~q ),
	.mem_66_0(\state_s1_agent_rsp_fifo|mem[0][66]~q ),
	.mem_65_0(\state_s1_agent_rsp_fifo|mem[0][65]~q ),
	.last_packet_beat1(\state_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(\state_s1_agent|uncompressor|last_packet_beat~2_combout ),
	.read(\state_s1_agent_rdata_fifo|read~0_combout ),
	.cp_ready1(\state_s1_agent|cp_ready~1_combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux cmd_mux(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.has_pending_responses(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.nxt_in_ready(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.Equal1(\router_001|Equal1~3_combout ),
	.last_channel_0(\hps_h2f_lw_axi_master_rd_limiter|last_channel[0]~q ),
	.src_valid(\cmd_mux|src_valid~0_combout ),
	.src_payload(\cmd_mux|src_payload~0_combout ),
	.src_payload1(\cmd_mux|src_payload~1_combout ),
	.src_payload2(\cmd_mux|src_payload~2_combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_demux_1 cmd_demux_001(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARADDR_16(h2f_lw_ARADDR_16),
	.h2f_lw_ARADDR_17(h2f_lw_ARADDR_17),
	.h2f_lw_ARADDR_18(h2f_lw_ARADDR_18),
	.nxt_in_ready(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.Equal5(\router_001|Equal5~0_combout ),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.nxt_in_ready3(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready4(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.sink_ready(\cmd_demux_001|sink_ready~0_combout ),
	.has_pending_responses(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_11(\cmd_mux_003|saved_grant[1]~q ),
	.Equal4(\router_001|Equal4~0_combout ),
	.Equal41(\router_001|Equal4~1_combout ),
	.nxt_in_ready5(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.sink_ready1(\cmd_demux_001|sink_ready~1_combout ),
	.nxt_in_ready6(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready7(\rbf_id_control_slave_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_12(\cmd_mux|saved_grant[1]~q ),
	.Equal12(\router_001|Equal1~2_combout ),
	.nxt_in_ready8(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready9(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_13(\cmd_mux_001|saved_grant[1]~q ),
	.WideOr01(\cmd_demux_001|WideOr0~0_combout ),
	.saved_grant_14(\cmd_mux_002|saved_grant[1]~q ),
	.Equal3(\router_001|Equal3~0_combout ),
	.nxt_in_ready10(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.sink_ready2(\cmd_demux_001|sink_ready~4_combout ),
	.saved_grant_15(\cmd_mux_004|saved_grant[1]~q ),
	.nxt_in_ready11(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.src_channel_4(\router_001|src_channel[4]~1_combout ),
	.sink_ready3(\cmd_demux_001|sink_ready~5_combout ),
	.WideOr02(\cmd_demux_001|WideOr0~combout ),
	.last_channel_3(\hps_h2f_lw_axi_master_rd_limiter|last_channel[3]~q ),
	.src3_valid(\cmd_demux_001|src3_valid~0_combout ),
	.src3_valid1(\cmd_demux_001|src3_valid~1_combout ),
	.last_channel_2(\hps_h2f_lw_axi_master_rd_limiter|last_channel[2]~q ),
	.src2_valid(\cmd_demux_001|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux_001|src2_valid~1_combout ),
	.last_channel_4(\hps_h2f_lw_axi_master_rd_limiter|last_channel[4]~q ),
	.src4_valid(\cmd_demux_001|src4_valid~0_combout ),
	.WideOr03(\cmd_demux_001|WideOr0~1_combout ),
	.src4_valid1(\cmd_demux_001|src4_valid~1_combout ));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_demux cmd_demux(
	.h2f_lw_AWVALID_0(h2f_lw_AWVALID_0),
	.h2f_lw_WVALID_0(h2f_lw_WVALID_0),
	.nxt_in_ready(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready1(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.nxt_in_ready2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready3(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready4(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.nxt_in_ready5(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal31(\router|Equal3~7_combout ),
	.Equal4(\router|Equal4~0_combout ),
	.has_pending_responses(\hps_h2f_lw_axi_master_wr_limiter|has_pending_responses~q ),
	.last_channel_2(\hps_h2f_lw_axi_master_wr_limiter|last_channel[2]~q ),
	.last_channel_4(\hps_h2f_lw_axi_master_wr_limiter|last_channel[4]~q ),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.saved_grant_01(\cmd_mux_002|saved_grant[0]~q ),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ),
	.saved_grant_02(\cmd_mux_004|saved_grant[0]~q ),
	.sink_ready2(\cmd_demux|sink_ready~2_combout ),
	.last_channel_3(\hps_h2f_lw_axi_master_wr_limiter|last_channel[3]~q ),
	.src3_valid(\cmd_demux|src3_valid~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src4_valid(\cmd_demux|src4_valid~0_combout ),
	.src4_valid1(\cmd_demux|src4_valid~1_combout ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ));

terminal_qsys_altera_merlin_burst_adapter_5 switches_s1_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.Add5(\hps_h2f_lw_axi_master_agent|Add5~9_sumout ),
	.Add51(\hps_h2f_lw_axi_master_agent|Add5~13_sumout ),
	.Equal5(\router_001|Equal5~0_combout ),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.mem_used_1(\switches_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_data_reg_60(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_narrow_reg(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.cp_ready(\switches_s1_agent|cp_ready~0_combout ),
	.nxt_in_ready(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.out_valid_reg(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.stateST_UNCOMP_WR_SUBBURST(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.nxt_out_eop(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.last_cycle(\cmd_mux_005|last_cycle~0_combout ),
	.Decoder1(\hps_h2f_lw_axi_master_agent|Decoder1~0_combout ),
	.out_byte_cnt_reg_2(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.cp_ready1(\switches_s1_agent|cp_ready~1_combout ),
	.out_uncomp_byte_cnt_reg_5(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_4(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_6(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_92(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.Selector10(\hps_h2f_lw_axi_master_agent|Selector10~0_combout ),
	.Selector101(\hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_34),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_24),
	.Add3(\hps_h2f_lw_axi_master_agent|Add3~3_combout ),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.Decoder11(\hps_h2f_lw_axi_master_agent|Decoder1~4_combout ),
	.src_payload(\cmd_mux_005|src_payload~0_combout ),
	.src_payload1(\cmd_mux_005|src_payload~1_combout ),
	.src_payload2(\cmd_mux_005|src_payload~2_combout ),
	.nxt_out_burstwrap_1(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[1]~0_combout ),
	.nxt_out_burstwrap_0(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_burst_adapter_2 leds_s1_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.nxt_in_ready(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.mem_used_1(\leds_s1_agent_rsp_fifo|mem_used[1]~q ),
	.in_narrow_reg(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_59(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.write(\leds_s1_agent_rsp_fifo|write~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.saved_grant_0(\cmd_mux_004|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.in_data_reg_0(in_data_reg_02),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_32),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_22),
	.in_data_reg_1(in_data_reg_112),
	.in_data_reg_2(in_data_reg_212),
	.in_data_reg_3(in_data_reg_33),
	.in_data_reg_4(in_data_reg_42),
	.in_data_reg_5(in_data_reg_52),
	.in_data_reg_6(in_data_reg_62),
	.in_data_reg_7(in_data_reg_72),
	.in_data_reg_8(in_data_reg_82),
	.in_data_reg_9(in_data_reg_92),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.write_cp_data_69(\hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.write_cp_data_68(\hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.write_cp_data_67(\hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.write_cp_data_66(\hps_h2f_lw_axi_master_agent|write_cp_data[66]~3_combout ),
	.write_cp_data_65(\hps_h2f_lw_axi_master_agent|write_cp_data[65]~4_combout ),
	.WideNor0(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.src_valid(\cmd_mux_004|src_valid~0_combout ),
	.src_valid1(\cmd_mux_004|src_valid~1_combout ),
	.src_payload_0(\cmd_mux_004|src_payload[0]~combout ),
	.nxt_out_eop(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready(\leds_s1_agent|cp_ready~0_combout ),
	.cp_ready1(\leds_s1_agent|cp_ready~1_combout ),
	.in_data_reg_60(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux_004|src_data[78]~combout ),
	.src_data_79(\cmd_mux_004|src_data[79]~combout ),
	.src_data_35(\cmd_mux_004|src_data[35]~combout ),
	.src_data_34(\cmd_mux_004|src_data[34]~combout ),
	.src_data_33(\cmd_mux_004|src_data[33]~combout ),
	.src_data_32(\cmd_mux_004|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_3(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_6(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.in_data_reg_92(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.base_address_3(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.base_address_2(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload(\cmd_mux_004|src_payload~0_combout ),
	.src_data_73(\cmd_mux_004|src_data[73]~combout ),
	.src_data_72(\cmd_mux_004|src_data[72]~combout ),
	.src_payload1(\cmd_mux_004|src_payload~1_combout ),
	.src_payload2(\cmd_mux_004|src_payload~2_combout ),
	.src_payload3(\cmd_mux_004|src_payload~3_combout ),
	.src_payload4(\cmd_mux_004|src_payload~4_combout ),
	.src_payload5(\cmd_mux_004|src_payload~5_combout ),
	.src_payload6(\cmd_mux_004|src_payload~6_combout ),
	.src_payload7(\cmd_mux_004|src_payload~7_combout ),
	.src_payload8(\cmd_mux_004|src_payload~8_combout ),
	.src_payload9(\cmd_mux_004|src_payload~9_combout ),
	.nxt_in_ready2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src_data_92(\cmd_mux_004|src_data[92]~combout ),
	.src_data_93(\cmd_mux_004|src_data[93]~combout ),
	.src_data_94(\cmd_mux_004|src_data[94]~combout ),
	.src_data_95(\cmd_mux_004|src_data[95]~combout ),
	.src_data_96(\cmd_mux_004|src_data[96]~combout ),
	.src_data_97(\cmd_mux_004|src_data[97]~combout ),
	.src_data_98(\cmd_mux_004|src_data[98]~combout ),
	.src_data_99(\cmd_mux_004|src_data[99]~combout ),
	.src_data_100(\cmd_mux_004|src_data[100]~combout ),
	.src_data_101(\cmd_mux_004|src_data[101]~combout ),
	.src_data_102(\cmd_mux_004|src_data[102]~combout ),
	.src_data_103(\cmd_mux_004|src_data[103]~combout ),
	.src_data_77(\cmd_mux_004|src_data[77]~combout ),
	.out_data_1(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~15_combout ),
	.src_data_71(\cmd_mux_004|src_data[71]~combout ),
	.out_data_0(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~16_combout ),
	.src_data_70(\cmd_mux_004|src_data[70]~combout ),
	.clk_clk(clk_clk));

terminal_qsys_altera_merlin_burst_adapter base_address_ddr_s1_burst_adapter(
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.nxt_in_ready(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.stateST_COMP_TRANS(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_COMP_TRANS~q ),
	.out_valid_reg(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_valid_reg~q ),
	.in_ready_hold(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.in_narrow_reg(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_narrow_reg~q ),
	.in_byteen_reg_3(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[3]~q ),
	.in_byteen_reg_2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[2]~q ),
	.in_byteen_reg_1(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[1]~q ),
	.in_byteen_reg_0(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_byteen_reg[0]~q ),
	.in_data_reg_59(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[59]~q ),
	.write(\base_address_ddr_s1_agent_rsp_fifo|write~0_combout ),
	.stateST_UNCOMP_WR_SUBBURST(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|state.ST_UNCOMP_WR_SUBBURST~q ),
	.nxt_in_ready1(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal4(\router|Equal4~0_combout ),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.in_data_reg_0(in_data_reg_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.Add2(\hps_h2f_lw_axi_master_agent|Add2~0_combout ),
	.Add21(\hps_h2f_lw_axi_master_agent|Add2~1_combout ),
	.Add22(\hps_h2f_lw_axi_master_agent|Add2~2_combout ),
	.src3_valid(\cmd_demux|src3_valid~0_combout ),
	.src_valid(\cmd_mux_003|src_valid~0_combout ),
	.src_payload_0(\cmd_mux_003|src_payload[0]~combout ),
	.nxt_out_eop(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_eop~0_combout ),
	.cp_ready(\base_address_ddr_s1_agent|cp_ready~2_combout ),
	.in_data_reg_60(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[60]~q ),
	.src_data_78(\cmd_mux_003|src_data[78]~combout ),
	.src_data_79(\cmd_mux_003|src_data[79]~combout ),
	.src_data_35(\cmd_mux_003|src_data[35]~combout ),
	.src_data_34(\cmd_mux_003|src_data[34]~combout ),
	.src_data_33(\cmd_mux_003|src_data[33]~combout ),
	.src_data_32(\cmd_mux_003|src_data[32]~combout ),
	.out_byte_cnt_reg_2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_4(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[4]~q ),
	.out_uncomp_byte_cnt_reg_3(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[3]~q ),
	.out_uncomp_byte_cnt_reg_2(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[2]~q ),
	.out_uncomp_byte_cnt_reg_5(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[5]~q ),
	.out_uncomp_byte_cnt_reg_6(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|out_uncomp_byte_cnt_reg[6]~q ),
	.write_cp_data_69(\hps_h2f_lw_axi_master_agent|write_cp_data[69]~0_combout ),
	.write_cp_data_68(\hps_h2f_lw_axi_master_agent|write_cp_data[68]~1_combout ),
	.write_cp_data_67(\hps_h2f_lw_axi_master_agent|write_cp_data[67]~2_combout ),
	.write_cp_data_66(\hps_h2f_lw_axi_master_agent|write_cp_data[66]~3_combout ),
	.write_cp_data_65(\hps_h2f_lw_axi_master_agent|write_cp_data[65]~4_combout ),
	.WideNor0(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|WideNor0~0_combout ),
	.in_data_reg_92(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[92]~q ),
	.in_data_reg_93(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[93]~q ),
	.in_data_reg_94(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[94]~q ),
	.in_data_reg_95(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[95]~q ),
	.in_data_reg_96(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[96]~q ),
	.in_data_reg_97(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[97]~q ),
	.in_data_reg_98(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[98]~q ),
	.in_data_reg_99(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[99]~q ),
	.in_data_reg_100(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[100]~q ),
	.in_data_reg_101(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[101]~q ),
	.in_data_reg_102(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[102]~q ),
	.in_data_reg_103(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_data_reg[103]~q ),
	.src_payload(\cmd_mux_003|src_payload~0_combout ),
	.src_data_73(\cmd_mux_003|src_data[73]~combout ),
	.base_address_3(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[3]~0_combout ),
	.src_data_72(\cmd_mux_003|src_data[72]~combout ),
	.base_address_2(\hps_h2f_lw_axi_master_agent|align_address_to_size|base_address[2]~1_combout ),
	.src_payload1(\cmd_mux_003|src_payload~1_combout ),
	.src_payload2(\cmd_mux_003|src_payload~2_combout ),
	.src_payload3(\cmd_mux_003|src_payload~3_combout ),
	.src_payload4(\cmd_mux_003|src_payload~4_combout ),
	.src_payload5(\cmd_mux_003|src_payload~5_combout ),
	.src_payload6(\cmd_mux_003|src_payload~6_combout ),
	.src_payload7(\cmd_mux_003|src_payload~7_combout ),
	.src_payload8(\cmd_mux_003|src_payload~8_combout ),
	.src_payload9(\cmd_mux_003|src_payload~9_combout ),
	.src_payload10(\cmd_mux_003|src_payload~10_combout ),
	.src_payload11(\cmd_mux_003|src_payload~11_combout ),
	.src_payload12(\cmd_mux_003|src_payload~12_combout ),
	.src_payload13(\cmd_mux_003|src_payload~13_combout ),
	.src_payload14(\cmd_mux_003|src_payload~14_combout ),
	.src_payload15(\cmd_mux_003|src_payload~15_combout ),
	.src_payload16(\cmd_mux_003|src_payload~16_combout ),
	.src_payload17(\cmd_mux_003|src_payload~17_combout ),
	.src_payload18(\cmd_mux_003|src_payload~18_combout ),
	.src_payload19(\cmd_mux_003|src_payload~19_combout ),
	.src_payload20(\cmd_mux_003|src_payload~20_combout ),
	.src_payload21(\cmd_mux_003|src_payload~21_combout ),
	.src_payload22(\cmd_mux_003|src_payload~22_combout ),
	.src_payload23(\cmd_mux_003|src_payload~23_combout ),
	.src_payload24(\cmd_mux_003|src_payload~24_combout ),
	.src_payload25(\cmd_mux_003|src_payload~25_combout ),
	.src_payload26(\cmd_mux_003|src_payload~26_combout ),
	.src_payload27(\cmd_mux_003|src_payload~27_combout ),
	.src_payload28(\cmd_mux_003|src_payload~28_combout ),
	.src_payload29(\cmd_mux_003|src_payload~29_combout ),
	.src_payload30(\cmd_mux_003|src_payload~30_combout ),
	.src_payload31(\cmd_mux_003|src_payload~31_combout ),
	.src_data_92(\cmd_mux_003|src_data[92]~combout ),
	.src_data_93(\cmd_mux_003|src_data[93]~combout ),
	.src_data_94(\cmd_mux_003|src_data[94]~combout ),
	.src_data_95(\cmd_mux_003|src_data[95]~combout ),
	.src_data_96(\cmd_mux_003|src_data[96]~combout ),
	.src_data_97(\cmd_mux_003|src_data[97]~combout ),
	.src_data_98(\cmd_mux_003|src_data[98]~combout ),
	.src_data_99(\cmd_mux_003|src_data[99]~combout ),
	.src_data_100(\cmd_mux_003|src_data[100]~combout ),
	.src_data_101(\cmd_mux_003|src_data[101]~combout ),
	.src_data_102(\cmd_mux_003|src_data[102]~combout ),
	.src_data_103(\cmd_mux_003|src_data[103]~combout ),
	.src_data_77(\cmd_mux_003|src_data[77]~combout ),
	.src_data_71(\cmd_mux_003|src_data[71]~combout ),
	.out_data_1(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[1]~15_combout ),
	.out_data_0(\hps_h2f_lw_axi_master_agent|align_address_to_size|out_data[0]~16_combout ),
	.src_data_70(\cmd_mux_003|src_data[70]~combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_mux_1 rsp_mux_001(
	.in_ready_hold(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|in_ready_hold~q ),
	.mem_57_0(\control_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_57_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_57_02(\leds_s1_agent_rsp_fifo|mem[0][57]~q ),
	.comb(\control_s1_agent|comb~0_combout ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.mem_117_0(\control_s1_agent_rsp_fifo|mem[0][117]~q ),
	.last_packet_beat(\control_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat1(\control_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb1(\base_address_ddr_s1_agent|comb~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.mem_117_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][117]~q ),
	.last_packet_beat2(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat3(\base_address_ddr_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.comb2(\leds_s1_agent|comb~0_combout ),
	.src1_valid2(\rsp_demux_004|src1_valid~0_combout ),
	.mem_117_02(\leds_s1_agent_rsp_fifo|mem[0][117]~q ),
	.last_packet_beat4(\leds_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat5(\leds_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_117_03(\switches_s1_agent_rsp_fifo|mem[0][117]~q ),
	.read_latency_shift_reg_0(\switches_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\switches_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty(\switches_s1_agent_rdata_fifo|empty~combout ),
	.mem_57_03(\switches_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_01(\switches_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat6(\switches_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat7(\switches_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_117_04(\state_s1_agent_rsp_fifo|mem[0][117]~q ),
	.read_latency_shift_reg_01(\state_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_02(\state_s1_agent_rdata_fifo|mem_used[0]~q ),
	.empty1(\state_s1_agent_rdata_fifo|empty~combout ),
	.mem_57_04(\state_s1_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_03(\state_s1_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat8(\state_s1_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat9(\state_s1_agent|uncompressor|last_packet_beat~1_combout ),
	.mem_117_05(\rbf_id_control_slave_agent_rsp_fifo|mem[0][117]~q ),
	.read_latency_shift_reg_02(\rbf_id_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_04(\rbf_id_control_slave_agent_rdata_fifo|mem_used[0]~q ),
	.empty2(\rbf_id_control_slave_agent_rdata_fifo|empty~combout ),
	.mem_57_05(\rbf_id_control_slave_agent_rsp_fifo|mem[0][57]~q ),
	.mem_used_05(\rbf_id_control_slave_agent_rsp_fifo|mem_used[0]~q ),
	.last_packet_beat10(\rbf_id_control_slave_agent|uncompressor|last_packet_beat~0_combout ),
	.last_packet_beat11(\rbf_id_control_slave_agent|uncompressor|last_packet_beat~1_combout ),
	.src_payload_0(src_payload_0),
	.WideOr11(WideOr11),
	.mem_92_0(\control_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_02(\leds_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_93_0(\control_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_02(\leds_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_94_0(\control_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_02(\leds_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_95_0(\control_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_02(\leds_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_96_0(\control_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_02(\leds_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_97_0(\control_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_02(\leds_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_98_0(\control_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_02(\leds_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_99_0(\control_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_02(\leds_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_100_0(\control_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_100_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_100_02(\leds_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_101_0(\control_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_02(\leds_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_102_0(\control_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_02(\leds_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_103_0(\control_s1_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_02(\leds_s1_agent_rsp_fifo|mem[0][103]~q ),
	.av_readdata_pre_0(\control_s1_translator|av_readdata_pre[0]~q ),
	.always4(\control_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_0(\control_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_01(\base_address_ddr_s1_translator|av_readdata_pre[0]~q ),
	.always41(\base_address_ddr_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_02(\leds_s1_translator|av_readdata_pre[0]~q ),
	.always42(\leds_s1_agent_rdata_fifo|always4~0_combout ),
	.mem_0_02(\leds_s1_agent_rdata_fifo|mem[0][0]~q ),
	.mem_0_03(\state_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_03(\state_s1_translator|av_readdata_pre[0]~q ),
	.mem_0_04(\switches_s1_agent_rdata_fifo|mem[0][0]~q ),
	.av_readdata_pre_04(\switches_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_1(\control_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_0(\control_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_11(\base_address_ddr_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_12(\leds_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_02(\leds_s1_agent_rdata_fifo|mem[0][1]~q ),
	.mem_1_03(\state_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_13(\state_s1_translator|av_readdata_pre[1]~q ),
	.mem_1_04(\switches_s1_agent_rdata_fifo|mem[0][1]~q ),
	.av_readdata_pre_14(\switches_s1_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_2(\control_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_0(\control_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_21(\base_address_ddr_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_22(\leds_s1_translator|av_readdata_pre[2]~q ),
	.mem_2_02(\leds_s1_agent_rdata_fifo|mem[0][2]~q ),
	.mem_2_03(\state_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_23(\state_s1_translator|av_readdata_pre[2]~q ),
	.mem_11_0(\rbf_id_control_slave_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_30(\rbf_id_control_slave_translator|av_readdata_pre[30]~q ),
	.mem_2_04(\switches_s1_agent_rdata_fifo|mem[0][2]~q ),
	.av_readdata_pre_24(\switches_s1_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_3(\control_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_0(\control_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_31(\base_address_ddr_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_32(\leds_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_02(\leds_s1_agent_rdata_fifo|mem[0][3]~q ),
	.mem_3_03(\state_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_33(\state_s1_translator|av_readdata_pre[3]~q ),
	.mem_3_04(\switches_s1_agent_rdata_fifo|mem[0][3]~q ),
	.av_readdata_pre_34(\switches_s1_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_4(\control_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_0(\control_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_41(\base_address_ddr_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_42(\leds_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_02(\leds_s1_agent_rdata_fifo|mem[0][4]~q ),
	.mem_4_03(\state_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_43(\state_s1_translator|av_readdata_pre[4]~q ),
	.mem_4_04(\switches_s1_agent_rdata_fifo|mem[0][4]~q ),
	.av_readdata_pre_44(\switches_s1_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_5(\control_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_0(\control_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_51(\base_address_ddr_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_52(\leds_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_02(\leds_s1_agent_rdata_fifo|mem[0][5]~q ),
	.mem_5_03(\state_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_53(\state_s1_translator|av_readdata_pre[5]~q ),
	.mem_5_04(\switches_s1_agent_rdata_fifo|mem[0][5]~q ),
	.av_readdata_pre_54(\switches_s1_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_6(\control_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_0(\control_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_61(\base_address_ddr_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_62(\leds_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_02(\leds_s1_agent_rdata_fifo|mem[0][6]~q ),
	.mem_6_03(\state_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_63(\state_s1_translator|av_readdata_pre[6]~q ),
	.mem_6_04(\switches_s1_agent_rdata_fifo|mem[0][6]~q ),
	.av_readdata_pre_64(\switches_s1_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_7(\control_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_0(\control_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_71(\base_address_ddr_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_72(\leds_s1_translator|av_readdata_pre[7]~q ),
	.mem_7_02(\leds_s1_agent_rdata_fifo|mem[0][7]~q ),
	.mem_7_03(\state_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_73(\state_s1_translator|av_readdata_pre[7]~q ),
	.mem_10_0(\rbf_id_control_slave_agent_rdata_fifo|mem[0][10]~q ),
	.mem_7_04(\switches_s1_agent_rdata_fifo|mem[0][7]~q ),
	.av_readdata_pre_74(\switches_s1_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_8(\control_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_0(\control_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_81(\base_address_ddr_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_82(\leds_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_02(\leds_s1_agent_rdata_fifo|mem[0][8]~q ),
	.mem_8_03(\state_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_83(\state_s1_translator|av_readdata_pre[8]~q ),
	.mem_8_04(\switches_s1_agent_rdata_fifo|mem[0][8]~q ),
	.av_readdata_pre_84(\switches_s1_translator|av_readdata_pre[8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_9(\state_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_91(\control_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_0(\control_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_92(\base_address_ddr_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_93(\leds_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_02(\leds_s1_agent_rdata_fifo|mem[0][9]~q ),
	.mem_9_03(\switches_s1_agent_rdata_fifo|mem[0][9]~q ),
	.av_readdata_pre_94(\switches_s1_translator|av_readdata_pre[9]~q ),
	.mem_9_04(\state_s1_agent_rdata_fifo|mem[0][9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_10(\control_s1_translator|av_readdata_pre[10]~q ),
	.mem_10_01(\control_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_101(\base_address_ddr_s1_translator|av_readdata_pre[10]~q ),
	.mem_10_02(\base_address_ddr_s1_agent_rdata_fifo|mem[0][10]~q ),
	.mem_10_03(\state_s1_agent_rdata_fifo|mem[0][10]~q ),
	.av_readdata_pre_102(\state_s1_translator|av_readdata_pre[10]~q ),
	.src_payload(src_payload12),
	.av_readdata_pre_111(\control_s1_translator|av_readdata_pre[11]~q ),
	.mem_11_01(\control_s1_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_112(\base_address_ddr_s1_translator|av_readdata_pre[11]~q ),
	.mem_11_02(\base_address_ddr_s1_agent_rdata_fifo|mem[0][11]~q ),
	.mem_11_03(\state_s1_agent_rdata_fifo|mem[0][11]~q ),
	.av_readdata_pre_113(\state_s1_translator|av_readdata_pre[11]~q ),
	.src_payload1(src_payload13),
	.av_readdata_pre_121(\base_address_ddr_s1_translator|av_readdata_pre[12]~q ),
	.mem_12_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_122(\control_s1_translator|av_readdata_pre[12]~q ),
	.mem_12_01(\control_s1_agent_rdata_fifo|mem[0][12]~q ),
	.mem_12_02(\state_s1_agent_rdata_fifo|mem[0][12]~q ),
	.av_readdata_pre_123(\state_s1_translator|av_readdata_pre[12]~q ),
	.src_payload2(src_payload14),
	.av_readdata_pre_131(\base_address_ddr_s1_translator|av_readdata_pre[13]~q ),
	.mem_13_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_132(\control_s1_translator|av_readdata_pre[13]~q ),
	.mem_13_01(\control_s1_agent_rdata_fifo|mem[0][13]~q ),
	.mem_13_02(\state_s1_agent_rdata_fifo|mem[0][13]~q ),
	.av_readdata_pre_133(\state_s1_translator|av_readdata_pre[13]~q ),
	.src_payload3(src_payload15),
	.av_readdata_pre_141(\base_address_ddr_s1_translator|av_readdata_pre[14]~q ),
	.mem_14_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_142(\control_s1_translator|av_readdata_pre[14]~q ),
	.mem_14_01(\control_s1_agent_rdata_fifo|mem[0][14]~q ),
	.mem_14_02(\state_s1_agent_rdata_fifo|mem[0][14]~q ),
	.av_readdata_pre_143(\state_s1_translator|av_readdata_pre[14]~q ),
	.src_payload4(src_payload16),
	.av_readdata_pre_15(\base_address_ddr_s1_translator|av_readdata_pre[15]~q ),
	.mem_15_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_151(\control_s1_translator|av_readdata_pre[15]~q ),
	.mem_15_01(\control_s1_agent_rdata_fifo|mem[0][15]~q ),
	.mem_15_02(\state_s1_agent_rdata_fifo|mem[0][15]~q ),
	.av_readdata_pre_152(\state_s1_translator|av_readdata_pre[15]~q ),
	.src_payload5(src_payload17),
	.av_readdata_pre_16(\base_address_ddr_s1_translator|av_readdata_pre[16]~q ),
	.mem_16_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_161(\control_s1_translator|av_readdata_pre[16]~q ),
	.mem_16_01(\control_s1_agent_rdata_fifo|mem[0][16]~q ),
	.mem_16_02(\state_s1_agent_rdata_fifo|mem[0][16]~q ),
	.av_readdata_pre_162(\state_s1_translator|av_readdata_pre[16]~q ),
	.src_payload6(src_payload18),
	.av_readdata_pre_17(\base_address_ddr_s1_translator|av_readdata_pre[17]~q ),
	.mem_17_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_171(\control_s1_translator|av_readdata_pre[17]~q ),
	.mem_17_01(\control_s1_agent_rdata_fifo|mem[0][17]~q ),
	.mem_17_02(\state_s1_agent_rdata_fifo|mem[0][17]~q ),
	.av_readdata_pre_172(\state_s1_translator|av_readdata_pre[17]~q ),
	.src_payload7(src_payload19),
	.av_readdata_pre_18(\base_address_ddr_s1_translator|av_readdata_pre[18]~q ),
	.mem_18_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_181(\control_s1_translator|av_readdata_pre[18]~q ),
	.mem_18_01(\control_s1_agent_rdata_fifo|mem[0][18]~q ),
	.mem_18_02(\state_s1_agent_rdata_fifo|mem[0][18]~q ),
	.av_readdata_pre_182(\state_s1_translator|av_readdata_pre[18]~q ),
	.src_payload8(src_payload20),
	.av_readdata_pre_19(\control_s1_translator|av_readdata_pre[19]~q ),
	.mem_19_0(\control_s1_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_191(\base_address_ddr_s1_translator|av_readdata_pre[19]~q ),
	.mem_19_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][19]~q ),
	.mem_19_02(\state_s1_agent_rdata_fifo|mem[0][19]~q ),
	.av_readdata_pre_192(\state_s1_translator|av_readdata_pre[19]~q ),
	.src_payload9(src_payload21),
	.av_readdata_pre_20(\control_s1_translator|av_readdata_pre[20]~q ),
	.mem_20_0(\control_s1_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_201(\base_address_ddr_s1_translator|av_readdata_pre[20]~q ),
	.mem_20_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][20]~q ),
	.mem_20_02(\state_s1_agent_rdata_fifo|mem[0][20]~q ),
	.av_readdata_pre_202(\state_s1_translator|av_readdata_pre[20]~q ),
	.src_payload10(src_payload22),
	.av_readdata_pre_211(\control_s1_translator|av_readdata_pre[21]~q ),
	.mem_21_0(\control_s1_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_212(\base_address_ddr_s1_translator|av_readdata_pre[21]~q ),
	.mem_21_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][21]~q ),
	.mem_21_02(\state_s1_agent_rdata_fifo|mem[0][21]~q ),
	.av_readdata_pre_213(\state_s1_translator|av_readdata_pre[21]~q ),
	.src_payload11(src_payload23),
	.av_readdata_pre_221(\base_address_ddr_s1_translator|av_readdata_pre[22]~q ),
	.mem_22_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_222(\control_s1_translator|av_readdata_pre[22]~q ),
	.mem_22_01(\control_s1_agent_rdata_fifo|mem[0][22]~q ),
	.mem_22_02(\state_s1_agent_rdata_fifo|mem[0][22]~q ),
	.av_readdata_pre_223(\state_s1_translator|av_readdata_pre[22]~q ),
	.src_payload12(src_payload24),
	.av_readdata_pre_231(\base_address_ddr_s1_translator|av_readdata_pre[23]~q ),
	.mem_23_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_232(\control_s1_translator|av_readdata_pre[23]~q ),
	.mem_23_01(\control_s1_agent_rdata_fifo|mem[0][23]~q ),
	.mem_23_02(\state_s1_agent_rdata_fifo|mem[0][23]~q ),
	.av_readdata_pre_233(\state_s1_translator|av_readdata_pre[23]~q ),
	.src_payload13(src_payload25),
	.av_readdata_pre_241(\control_s1_translator|av_readdata_pre[24]~q ),
	.mem_24_0(\control_s1_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_242(\base_address_ddr_s1_translator|av_readdata_pre[24]~q ),
	.mem_24_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][24]~q ),
	.mem_24_02(\state_s1_agent_rdata_fifo|mem[0][24]~q ),
	.av_readdata_pre_243(\state_s1_translator|av_readdata_pre[24]~q ),
	.src_payload14(src_payload26),
	.av_readdata_pre_25(\base_address_ddr_s1_translator|av_readdata_pre[25]~q ),
	.mem_25_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_251(\control_s1_translator|av_readdata_pre[25]~q ),
	.mem_25_01(\control_s1_agent_rdata_fifo|mem[0][25]~q ),
	.mem_25_02(\state_s1_agent_rdata_fifo|mem[0][25]~q ),
	.av_readdata_pre_252(\state_s1_translator|av_readdata_pre[25]~q ),
	.src_payload15(src_payload27),
	.av_readdata_pre_26(\base_address_ddr_s1_translator|av_readdata_pre[26]~q ),
	.mem_26_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_261(\control_s1_translator|av_readdata_pre[26]~q ),
	.mem_26_01(\control_s1_agent_rdata_fifo|mem[0][26]~q ),
	.mem_26_02(\state_s1_agent_rdata_fifo|mem[0][26]~q ),
	.av_readdata_pre_262(\state_s1_translator|av_readdata_pre[26]~q ),
	.src_payload16(src_payload28),
	.av_readdata_pre_27(\control_s1_translator|av_readdata_pre[27]~q ),
	.mem_27_0(\control_s1_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_271(\base_address_ddr_s1_translator|av_readdata_pre[27]~q ),
	.mem_27_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][27]~q ),
	.mem_27_02(\state_s1_agent_rdata_fifo|mem[0][27]~q ),
	.av_readdata_pre_272(\state_s1_translator|av_readdata_pre[27]~q ),
	.src_payload17(src_payload29),
	.av_readdata_pre_28(\control_s1_translator|av_readdata_pre[28]~q ),
	.mem_28_0(\control_s1_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_281(\base_address_ddr_s1_translator|av_readdata_pre[28]~q ),
	.mem_28_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][28]~q ),
	.mem_28_02(\state_s1_agent_rdata_fifo|mem[0][28]~q ),
	.av_readdata_pre_282(\state_s1_translator|av_readdata_pre[28]~q ),
	.src_payload18(src_payload30),
	.av_readdata_pre_29(\base_address_ddr_s1_translator|av_readdata_pre[29]~q ),
	.mem_29_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_291(\control_s1_translator|av_readdata_pre[29]~q ),
	.mem_29_01(\control_s1_agent_rdata_fifo|mem[0][29]~q ),
	.mem_29_02(\state_s1_agent_rdata_fifo|mem[0][29]~q ),
	.av_readdata_pre_292(\state_s1_translator|av_readdata_pre[29]~q ),
	.src_payload19(src_payload31),
	.av_readdata_pre_301(\control_s1_translator|av_readdata_pre[30]~q ),
	.mem_30_0(\control_s1_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_302(\base_address_ddr_s1_translator|av_readdata_pre[30]~q ),
	.mem_30_01(\base_address_ddr_s1_agent_rdata_fifo|mem[0][30]~q ),
	.mem_30_02(\state_s1_agent_rdata_fifo|mem[0][30]~q ),
	.av_readdata_pre_303(\state_s1_translator|av_readdata_pre[30]~q ),
	.src_payload20(src_payload32),
	.av_readdata_pre_311(\base_address_ddr_s1_translator|av_readdata_pre[31]~q ),
	.mem_31_0(\base_address_ddr_s1_agent_rdata_fifo|mem[0][31]~q ),
	.av_readdata_pre_312(\control_s1_translator|av_readdata_pre[31]~q ),
	.mem_31_01(\control_s1_agent_rdata_fifo|mem[0][31]~q ),
	.mem_31_02(\state_s1_agent_rdata_fifo|mem[0][31]~q ),
	.av_readdata_pre_313(\state_s1_translator|av_readdata_pre[31]~q ),
	.src_payload21(src_payload33),
	.mem_92_03(\switches_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_05(\state_s1_agent_rsp_fifo|mem[0][92]~q ),
	.src_data_92(src_data_92),
	.mem_93_03(\switches_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_05(\state_s1_agent_rsp_fifo|mem[0][93]~q ),
	.src_data_93(src_data_93),
	.mem_94_03(\switches_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_05(\state_s1_agent_rsp_fifo|mem[0][94]~q ),
	.src_data_94(src_data_94),
	.mem_95_03(\switches_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_05(\state_s1_agent_rsp_fifo|mem[0][95]~q ),
	.src_data_95(src_data_95),
	.mem_96_03(\switches_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_05(\state_s1_agent_rsp_fifo|mem[0][96]~q ),
	.src_data_96(src_data_96),
	.mem_97_03(\switches_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_05(\state_s1_agent_rsp_fifo|mem[0][97]~q ),
	.src_data_97(src_data_97),
	.mem_98_03(\switches_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_05(\state_s1_agent_rsp_fifo|mem[0][98]~q ),
	.src_data_98(src_data_98),
	.mem_99_03(\switches_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_05(\state_s1_agent_rsp_fifo|mem[0][99]~q ),
	.src_data_99(src_data_99),
	.mem_100_03(\switches_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_100_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][100]~q ),
	.mem_100_05(\state_s1_agent_rsp_fifo|mem[0][100]~q ),
	.src_data_100(src_data_100),
	.mem_101_03(\switches_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_05(\state_s1_agent_rsp_fifo|mem[0][101]~q ),
	.src_data_101(src_data_101),
	.mem_102_03(\switches_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_05(\state_s1_agent_rsp_fifo|mem[0][102]~q ),
	.src_data_102(src_data_102),
	.mem_103_03(\switches_s1_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_04(\rbf_id_control_slave_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_05(\state_s1_agent_rsp_fifo|mem[0][103]~q ),
	.src_data_103(src_data_103),
	.src_payload22(\rsp_mux_001|src_payload~75_combout ));

terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_mux rsp_mux(
	.src0_valid(\rsp_demux_002|src0_valid~combout ),
	.src0_valid1(\rsp_demux_003|src0_valid~combout ),
	.src0_valid2(\rsp_demux_004|src0_valid~combout ),
	.WideOr11(WideOr1),
	.mem_92_0(\control_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][92]~q ),
	.mem_92_02(\leds_s1_agent_rsp_fifo|mem[0][92]~q ),
	.src_payload(src_payload),
	.mem_93_0(\control_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][93]~q ),
	.mem_93_02(\leds_s1_agent_rsp_fifo|mem[0][93]~q ),
	.src_payload1(src_payload1),
	.mem_94_0(\control_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][94]~q ),
	.mem_94_02(\leds_s1_agent_rsp_fifo|mem[0][94]~q ),
	.src_payload2(src_payload2),
	.mem_95_0(\control_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][95]~q ),
	.mem_95_02(\leds_s1_agent_rsp_fifo|mem[0][95]~q ),
	.src_payload3(src_payload3),
	.mem_96_0(\control_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][96]~q ),
	.mem_96_02(\leds_s1_agent_rsp_fifo|mem[0][96]~q ),
	.src_payload4(src_payload4),
	.mem_97_0(\control_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][97]~q ),
	.mem_97_02(\leds_s1_agent_rsp_fifo|mem[0][97]~q ),
	.src_payload5(src_payload5),
	.mem_98_0(\control_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][98]~q ),
	.mem_98_02(\leds_s1_agent_rsp_fifo|mem[0][98]~q ),
	.src_payload6(src_payload6),
	.mem_99_0(\control_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][99]~q ),
	.mem_99_02(\leds_s1_agent_rsp_fifo|mem[0][99]~q ),
	.src_payload7(src_payload7),
	.mem_100_0(\control_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_100_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][100]~q ),
	.mem_100_02(\leds_s1_agent_rsp_fifo|mem[0][100]~q ),
	.src_payload8(src_payload8),
	.mem_101_0(\control_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][101]~q ),
	.mem_101_02(\leds_s1_agent_rsp_fifo|mem[0][101]~q ),
	.src_payload9(src_payload9),
	.mem_102_0(\control_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][102]~q ),
	.mem_102_02(\leds_s1_agent_rsp_fifo|mem[0][102]~q ),
	.src_payload10(src_payload10),
	.mem_103_0(\control_s1_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_01(\base_address_ddr_s1_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_02(\leds_s1_agent_rsp_fifo|mem[0][103]~q ),
	.src_payload11(src_payload11));

terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_demux_4 rsp_demux_004(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\leds_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\leds_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\leds_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\leds_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\leds_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\leds_s1_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux_004|src0_valid~combout ),
	.src1_valid(\rsp_demux_004|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_004|WideOr0~0_combout ));

terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_demux_3 rsp_demux_003(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\base_address_ddr_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\base_address_ddr_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\base_address_ddr_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\base_address_ddr_s1_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux_003|src0_valid~combout ),
	.src1_valid(\rsp_demux_003|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_003|WideOr0~0_combout ));

terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_demux_2 rsp_demux_002(
	.h2f_lw_BREADY_0(h2f_lw_BREADY_0),
	.h2f_lw_RREADY_0(h2f_lw_RREADY_0),
	.read_latency_shift_reg_0(\control_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_0(\control_s1_agent_rdata_fifo|mem_used[0]~q ),
	.mem_116_0(\control_s1_agent_rsp_fifo|mem[0][116]~q ),
	.mem_used_01(\control_s1_agent_rsp_fifo|mem_used[0]~q ),
	.mem_59_0(\control_s1_agent_rsp_fifo|mem[0][59]~q ),
	.mem_57_0(\control_s1_agent_rsp_fifo|mem[0][57]~q ),
	.src0_valid1(\rsp_demux_002|src0_valid~combout ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.WideOr0(\rsp_demux_002|WideOr0~0_combout ));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_5 cmd_mux_005(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.Equal5(\router_001|Equal5~0_combout ),
	.saved_grant_1(\cmd_mux_005|saved_grant[1]~q ),
	.nxt_in_ready(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.has_pending_responses(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.last_channel_5(\hps_h2f_lw_axi_master_rd_limiter|last_channel[5]~q ),
	.last_cycle(\cmd_mux_005|last_cycle~0_combout ),
	.src_payload(\cmd_mux_005|src_payload~0_combout ),
	.src_payload1(\cmd_mux_005|src_payload~1_combout ),
	.src_payload2(\cmd_mux_005|src_payload~2_combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_4 cmd_mux_004(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.nxt_in_ready(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.has_pending_responses(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.saved_grant_1(\cmd_mux_004|saved_grant[1]~q ),
	.nxt_in_ready1(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.src_channel_4(\router_001|src_channel[4]~1_combout ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal31(\router|Equal3~7_combout ),
	.Equal4(\router|Equal4~0_combout ),
	.saved_grant_0(\cmd_mux_004|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.src4_valid(\cmd_demux|src4_valid~0_combout ),
	.src4_valid1(\cmd_demux|src4_valid~1_combout ),
	.last_channel_4(\hps_h2f_lw_axi_master_rd_limiter|last_channel[4]~q ),
	.src4_valid2(\cmd_demux_001|src4_valid~0_combout ),
	.src_valid(\cmd_mux_004|src_valid~0_combout ),
	.src_valid1(\cmd_mux_004|src_valid~1_combout ),
	.src_payload_0(\cmd_mux_004|src_payload[0]~combout ),
	.src_data_78(\cmd_mux_004|src_data[78]~combout ),
	.src_data_79(\cmd_mux_004|src_data[79]~combout ),
	.src_data_35(\cmd_mux_004|src_data[35]~combout ),
	.src_data_34(\cmd_mux_004|src_data[34]~combout ),
	.src_data_33(\cmd_mux_004|src_data[33]~combout ),
	.src_data_32(\cmd_mux_004|src_data[32]~combout ),
	.Selector3(\hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_h2f_lw_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_004|src_payload~0_combout ),
	.src_data_73(\cmd_mux_004|src_data[73]~combout ),
	.src_data_72(\cmd_mux_004|src_data[72]~combout ),
	.src_payload1(\cmd_mux_004|src_payload~1_combout ),
	.src_payload2(\cmd_mux_004|src_payload~2_combout ),
	.src_payload3(\cmd_mux_004|src_payload~3_combout ),
	.src_payload4(\cmd_mux_004|src_payload~4_combout ),
	.src_payload5(\cmd_mux_004|src_payload~5_combout ),
	.src_payload6(\cmd_mux_004|src_payload~6_combout ),
	.src_payload7(\cmd_mux_004|src_payload~7_combout ),
	.src_payload8(\cmd_mux_004|src_payload~8_combout ),
	.src_payload9(\cmd_mux_004|src_payload~9_combout ),
	.nxt_in_ready2(\leds_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.src4_valid3(\cmd_demux_001|src4_valid~1_combout ),
	.src_data_92(\cmd_mux_004|src_data[92]~combout ),
	.src_data_93(\cmd_mux_004|src_data[93]~combout ),
	.src_data_94(\cmd_mux_004|src_data[94]~combout ),
	.src_data_95(\cmd_mux_004|src_data[95]~combout ),
	.src_data_96(\cmd_mux_004|src_data[96]~combout ),
	.src_data_97(\cmd_mux_004|src_data[97]~combout ),
	.src_data_98(\cmd_mux_004|src_data[98]~combout ),
	.src_data_99(\cmd_mux_004|src_data[99]~combout ),
	.src_data_100(\cmd_mux_004|src_data[100]~combout ),
	.src_data_101(\cmd_mux_004|src_data[101]~combout ),
	.src_data_102(\cmd_mux_004|src_data[102]~combout ),
	.src_data_103(\cmd_mux_004|src_data[103]~combout ),
	.src_data_77(\cmd_mux_004|src_data[77]~combout ),
	.Selector5(\hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.src_data_71(\cmd_mux_004|src_data[71]~combout ),
	.Selector6(\hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.nxt_out_burstwrap_0(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ),
	.src_data_70(\cmd_mux_004|src_data[70]~combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_3 cmd_mux_003(
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_ARADDR_16(h2f_lw_ARADDR_16),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.nxt_in_ready(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.saved_grant_1(\cmd_mux_003|saved_grant[1]~q ),
	.Equal4(\router_001|Equal4~0_combout ),
	.nxt_in_ready1(\base_address_ddr_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal41(\router|Equal4~0_combout ),
	.saved_grant_0(\cmd_mux_003|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src3_valid(\cmd_demux|src3_valid~0_combout ),
	.src3_valid1(\cmd_demux_001|src3_valid~0_combout ),
	.src3_valid2(\cmd_demux_001|src3_valid~1_combout ),
	.src_valid(\cmd_mux_003|src_valid~0_combout ),
	.src_payload_0(\cmd_mux_003|src_payload[0]~combout ),
	.src_data_78(\cmd_mux_003|src_data[78]~combout ),
	.src_data_79(\cmd_mux_003|src_data[79]~combout ),
	.src_data_35(\cmd_mux_003|src_data[35]~combout ),
	.src_data_34(\cmd_mux_003|src_data[34]~combout ),
	.src_data_33(\cmd_mux_003|src_data[33]~combout ),
	.src_data_32(\cmd_mux_003|src_data[32]~combout ),
	.src_payload(\cmd_mux_003|src_payload~0_combout ),
	.Selector3(\hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.src_data_73(\cmd_mux_003|src_data[73]~combout ),
	.Selector4(\hps_h2f_lw_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.src_data_72(\cmd_mux_003|src_data[72]~combout ),
	.src_payload1(\cmd_mux_003|src_payload~1_combout ),
	.src_payload2(\cmd_mux_003|src_payload~2_combout ),
	.src_payload3(\cmd_mux_003|src_payload~3_combout ),
	.src_payload4(\cmd_mux_003|src_payload~4_combout ),
	.src_payload5(\cmd_mux_003|src_payload~5_combout ),
	.src_payload6(\cmd_mux_003|src_payload~6_combout ),
	.src_payload7(\cmd_mux_003|src_payload~7_combout ),
	.src_payload8(\cmd_mux_003|src_payload~8_combout ),
	.src_payload9(\cmd_mux_003|src_payload~9_combout ),
	.src_payload10(\cmd_mux_003|src_payload~10_combout ),
	.src_payload11(\cmd_mux_003|src_payload~11_combout ),
	.src_payload12(\cmd_mux_003|src_payload~12_combout ),
	.src_payload13(\cmd_mux_003|src_payload~13_combout ),
	.src_payload14(\cmd_mux_003|src_payload~14_combout ),
	.src_payload15(\cmd_mux_003|src_payload~15_combout ),
	.src_payload16(\cmd_mux_003|src_payload~16_combout ),
	.src_payload17(\cmd_mux_003|src_payload~17_combout ),
	.src_payload18(\cmd_mux_003|src_payload~18_combout ),
	.src_payload19(\cmd_mux_003|src_payload~19_combout ),
	.src_payload20(\cmd_mux_003|src_payload~20_combout ),
	.src_payload21(\cmd_mux_003|src_payload~21_combout ),
	.src_payload22(\cmd_mux_003|src_payload~22_combout ),
	.src_payload23(\cmd_mux_003|src_payload~23_combout ),
	.src_payload24(\cmd_mux_003|src_payload~24_combout ),
	.src_payload25(\cmd_mux_003|src_payload~25_combout ),
	.src_payload26(\cmd_mux_003|src_payload~26_combout ),
	.src_payload27(\cmd_mux_003|src_payload~27_combout ),
	.src_payload28(\cmd_mux_003|src_payload~28_combout ),
	.src_payload29(\cmd_mux_003|src_payload~29_combout ),
	.src_payload30(\cmd_mux_003|src_payload~30_combout ),
	.src_payload31(\cmd_mux_003|src_payload~31_combout ),
	.src_data_92(\cmd_mux_003|src_data[92]~combout ),
	.src_data_93(\cmd_mux_003|src_data[93]~combout ),
	.src_data_94(\cmd_mux_003|src_data[94]~combout ),
	.src_data_95(\cmd_mux_003|src_data[95]~combout ),
	.src_data_96(\cmd_mux_003|src_data[96]~combout ),
	.src_data_97(\cmd_mux_003|src_data[97]~combout ),
	.src_data_98(\cmd_mux_003|src_data[98]~combout ),
	.src_data_99(\cmd_mux_003|src_data[99]~combout ),
	.src_data_100(\cmd_mux_003|src_data[100]~combout ),
	.src_data_101(\cmd_mux_003|src_data[101]~combout ),
	.src_data_102(\cmd_mux_003|src_data[102]~combout ),
	.src_data_103(\cmd_mux_003|src_data[103]~combout ),
	.src_data_77(\cmd_mux_003|src_data[77]~combout ),
	.Selector5(\hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.src_data_71(\cmd_mux_003|src_data[71]~combout ),
	.Selector6(\hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.nxt_out_burstwrap_0(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ),
	.src_data_70(\cmd_mux_003|src_data[70]~combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_2 cmd_mux_002(
	.h2f_lw_WLAST_0(h2f_lw_WLAST_0),
	.h2f_lw_ARADDR_17(h2f_lw_ARADDR_17),
	.h2f_lw_ARID_0(h2f_lw_ARID_0),
	.h2f_lw_ARID_1(h2f_lw_ARID_1),
	.h2f_lw_ARID_2(h2f_lw_ARID_2),
	.h2f_lw_ARID_3(h2f_lw_ARID_3),
	.h2f_lw_ARID_4(h2f_lw_ARID_4),
	.h2f_lw_ARID_5(h2f_lw_ARID_5),
	.h2f_lw_ARID_6(h2f_lw_ARID_6),
	.h2f_lw_ARID_7(h2f_lw_ARID_7),
	.h2f_lw_ARID_8(h2f_lw_ARID_8),
	.h2f_lw_ARID_9(h2f_lw_ARID_9),
	.h2f_lw_ARID_10(h2f_lw_ARID_10),
	.h2f_lw_ARID_11(h2f_lw_ARID_11),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.h2f_lw_AWID_0(h2f_lw_AWID_0),
	.h2f_lw_AWID_1(h2f_lw_AWID_1),
	.h2f_lw_AWID_2(h2f_lw_AWID_2),
	.h2f_lw_AWID_3(h2f_lw_AWID_3),
	.h2f_lw_AWID_4(h2f_lw_AWID_4),
	.h2f_lw_AWID_5(h2f_lw_AWID_5),
	.h2f_lw_AWID_6(h2f_lw_AWID_6),
	.h2f_lw_AWID_7(h2f_lw_AWID_7),
	.h2f_lw_AWID_8(h2f_lw_AWID_8),
	.h2f_lw_AWID_9(h2f_lw_AWID_9),
	.h2f_lw_AWID_10(h2f_lw_AWID_10),
	.h2f_lw_AWID_11(h2f_lw_AWID_11),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.h2f_lw_WDATA_0(h2f_lw_WDATA_0),
	.h2f_lw_WDATA_1(h2f_lw_WDATA_1),
	.h2f_lw_WDATA_2(h2f_lw_WDATA_2),
	.h2f_lw_WDATA_3(h2f_lw_WDATA_3),
	.h2f_lw_WDATA_4(h2f_lw_WDATA_4),
	.h2f_lw_WDATA_5(h2f_lw_WDATA_5),
	.h2f_lw_WDATA_6(h2f_lw_WDATA_6),
	.h2f_lw_WDATA_7(h2f_lw_WDATA_7),
	.h2f_lw_WDATA_8(h2f_lw_WDATA_8),
	.h2f_lw_WDATA_9(h2f_lw_WDATA_9),
	.h2f_lw_WDATA_10(h2f_lw_WDATA_10),
	.h2f_lw_WDATA_11(h2f_lw_WDATA_11),
	.h2f_lw_WDATA_12(h2f_lw_WDATA_12),
	.h2f_lw_WDATA_13(h2f_lw_WDATA_13),
	.h2f_lw_WDATA_14(h2f_lw_WDATA_14),
	.h2f_lw_WDATA_15(h2f_lw_WDATA_15),
	.h2f_lw_WDATA_16(h2f_lw_WDATA_16),
	.h2f_lw_WDATA_17(h2f_lw_WDATA_17),
	.h2f_lw_WDATA_18(h2f_lw_WDATA_18),
	.h2f_lw_WDATA_19(h2f_lw_WDATA_19),
	.h2f_lw_WDATA_20(h2f_lw_WDATA_20),
	.h2f_lw_WDATA_21(h2f_lw_WDATA_21),
	.h2f_lw_WDATA_22(h2f_lw_WDATA_22),
	.h2f_lw_WDATA_23(h2f_lw_WDATA_23),
	.h2f_lw_WDATA_24(h2f_lw_WDATA_24),
	.h2f_lw_WDATA_25(h2f_lw_WDATA_25),
	.h2f_lw_WDATA_26(h2f_lw_WDATA_26),
	.h2f_lw_WDATA_27(h2f_lw_WDATA_27),
	.h2f_lw_WDATA_28(h2f_lw_WDATA_28),
	.h2f_lw_WDATA_29(h2f_lw_WDATA_29),
	.h2f_lw_WDATA_30(h2f_lw_WDATA_30),
	.h2f_lw_WDATA_31(h2f_lw_WDATA_31),
	.h2f_lw_WSTRB_0(h2f_lw_WSTRB_0),
	.h2f_lw_WSTRB_1(h2f_lw_WSTRB_1),
	.h2f_lw_WSTRB_2(h2f_lw_WSTRB_2),
	.h2f_lw_WSTRB_3(h2f_lw_WSTRB_3),
	.nxt_in_ready(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~2_combout ),
	.Equal1(\router_001|Equal1~0_combout ),
	.Equal11(\router_001|Equal1~1_combout ),
	.Equal12(\router_001|Equal1~2_combout ),
	.saved_grant_1(\cmd_mux_002|saved_grant[1]~q ),
	.nxt_in_ready1(\control_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.Equal3(\router|Equal3~6_combout ),
	.Equal31(\router|Equal3~7_combout ),
	.saved_grant_0(\cmd_mux_002|saved_grant[0]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out1),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux_001|src2_valid~0_combout ),
	.src2_valid2(\cmd_demux_001|src2_valid~1_combout ),
	.src_valid(\cmd_mux_002|src_valid~0_combout ),
	.src_payload_0(\cmd_mux_002|src_payload[0]~combout ),
	.src_data_78(\cmd_mux_002|src_data[78]~combout ),
	.src_data_79(\cmd_mux_002|src_data[79]~combout ),
	.src_data_35(\cmd_mux_002|src_data[35]~combout ),
	.src_data_34(\cmd_mux_002|src_data[34]~combout ),
	.src_data_33(\cmd_mux_002|src_data[33]~combout ),
	.src_data_32(\cmd_mux_002|src_data[32]~combout ),
	.Selector3(\hps_h2f_lw_axi_master_agent|Selector3~0_combout ),
	.Selector10(\hps_h2f_lw_axi_master_agent|Selector10~1_combout ),
	.Selector4(\hps_h2f_lw_axi_master_agent|Selector4~1_combout ),
	.Selector11(\hps_h2f_lw_axi_master_agent|Selector11~1_combout ),
	.src_payload(\cmd_mux_002|src_payload~0_combout ),
	.src_data_73(\cmd_mux_002|src_data[73]~combout ),
	.src_data_72(\cmd_mux_002|src_data[72]~combout ),
	.src_payload1(\cmd_mux_002|src_payload~1_combout ),
	.src_payload2(\cmd_mux_002|src_payload~2_combout ),
	.src_payload3(\cmd_mux_002|src_payload~3_combout ),
	.src_payload4(\cmd_mux_002|src_payload~4_combout ),
	.src_payload5(\cmd_mux_002|src_payload~5_combout ),
	.src_payload6(\cmd_mux_002|src_payload~6_combout ),
	.src_payload7(\cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\cmd_mux_002|src_payload~31_combout ),
	.src_data_92(\cmd_mux_002|src_data[92]~combout ),
	.src_data_93(\cmd_mux_002|src_data[93]~combout ),
	.src_data_94(\cmd_mux_002|src_data[94]~combout ),
	.src_data_95(\cmd_mux_002|src_data[95]~combout ),
	.src_data_96(\cmd_mux_002|src_data[96]~combout ),
	.src_data_97(\cmd_mux_002|src_data[97]~combout ),
	.src_data_98(\cmd_mux_002|src_data[98]~combout ),
	.src_data_99(\cmd_mux_002|src_data[99]~combout ),
	.src_data_100(\cmd_mux_002|src_data[100]~combout ),
	.src_data_101(\cmd_mux_002|src_data[101]~combout ),
	.src_data_102(\cmd_mux_002|src_data[102]~combout ),
	.src_data_103(\cmd_mux_002|src_data[103]~combout ),
	.src_data_77(\cmd_mux_002|src_data[77]~combout ),
	.Selector5(\hps_h2f_lw_axi_master_agent|Selector5~1_combout ),
	.Selector12(\hps_h2f_lw_axi_master_agent|Selector12~0_combout ),
	.src_data_71(\cmd_mux_002|src_data[71]~combout ),
	.Selector6(\hps_h2f_lw_axi_master_agent|Selector6~0_combout ),
	.nxt_out_burstwrap_0(\switches_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_out_burstwrap[0]~2_combout ),
	.src_data_70(\cmd_mux_002|src_data[70]~combout ),
	.clk_clk(clk_clk));

terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_1 cmd_mux_001(
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARSIZE_0(h2f_lw_ARSIZE_0),
	.h2f_lw_ARSIZE_1(h2f_lw_ARSIZE_1),
	.h2f_lw_ARSIZE_2(h2f_lw_ARSIZE_2),
	.has_pending_responses(\hps_h2f_lw_axi_master_rd_limiter|has_pending_responses~q ),
	.nxt_in_ready(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~0_combout ),
	.nxt_in_ready1(\state_s1_burst_adapter|altera_merlin_burst_adapter_13_1.burst_adapter|nxt_in_ready~1_combout ),
	.saved_grant_1(\cmd_mux_001|saved_grant[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal2(\router_001|Equal2~0_combout ),
	.last_channel_1(\hps_h2f_lw_axi_master_rd_limiter|last_channel[1]~q ),
	.src_valid(\cmd_mux_001|src_valid~0_combout ),
	.src_valid1(\cmd_mux_001|src_valid~1_combout ),
	.src_payload(\cmd_mux_001|src_payload~0_combout ),
	.src_payload1(\cmd_mux_001|src_payload~1_combout ),
	.src_payload2(\cmd_mux_001|src_payload~2_combout ),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_avalon_sc_fifo (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_9,
	mem_9_0,
	av_readdata_pre_10,
	mem_10_0,
	av_readdata_pre_11,
	mem_11_0,
	av_readdata_pre_12,
	mem_12_0,
	av_readdata_pre_13,
	mem_13_0,
	av_readdata_pre_14,
	mem_14_0,
	av_readdata_pre_15,
	mem_15_0,
	av_readdata_pre_16,
	mem_16_0,
	av_readdata_pre_17,
	mem_17_0,
	av_readdata_pre_18,
	mem_18_0,
	av_readdata_pre_19,
	mem_19_0,
	av_readdata_pre_20,
	mem_20_0,
	av_readdata_pre_21,
	mem_21_0,
	av_readdata_pre_22,
	mem_22_0,
	av_readdata_pre_23,
	mem_23_0,
	av_readdata_pre_24,
	mem_24_0,
	av_readdata_pre_25,
	mem_25_0,
	av_readdata_pre_26,
	mem_26_0,
	av_readdata_pre_27,
	mem_27_0,
	av_readdata_pre_28,
	mem_28_0,
	av_readdata_pre_29,
	mem_29_0,
	av_readdata_pre_30,
	mem_30_0,
	av_readdata_pre_31,
	mem_31_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	always4;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	av_readdata_pre_8;
output 	mem_8_0;
input 	av_readdata_pre_9;
output 	mem_9_0;
input 	av_readdata_pre_10;
output 	mem_10_0;
input 	av_readdata_pre_11;
output 	mem_11_0;
input 	av_readdata_pre_12;
output 	mem_12_0;
input 	av_readdata_pre_13;
output 	mem_13_0;
input 	av_readdata_pre_14;
output 	mem_14_0;
input 	av_readdata_pre_15;
output 	mem_15_0;
input 	av_readdata_pre_16;
output 	mem_16_0;
input 	av_readdata_pre_17;
output 	mem_17_0;
input 	av_readdata_pre_18;
output 	mem_18_0;
input 	av_readdata_pre_19;
output 	mem_19_0;
input 	av_readdata_pre_20;
output 	mem_20_0;
input 	av_readdata_pre_21;
output 	mem_21_0;
input 	av_readdata_pre_22;
output 	mem_22_0;
input 	av_readdata_pre_23;
output 	mem_23_0;
input 	av_readdata_pre_24;
output 	mem_24_0;
input 	av_readdata_pre_25;
output 	mem_25_0;
input 	av_readdata_pre_26;
output 	mem_26_0;
input 	av_readdata_pre_27;
output 	mem_27_0;
input 	av_readdata_pre_28;
output 	mem_28_0;
input 	av_readdata_pre_29;
output 	mem_29_0;
input 	av_readdata_pre_30;
output 	mem_30_0;
input 	av_readdata_pre_31;
output 	mem_31_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!av_readdata_pre_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!av_readdata_pre_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!av_readdata_pre_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!av_readdata_pre_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!av_readdata_pre_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!av_readdata_pre_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!av_readdata_pre_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!av_readdata_pre_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!av_readdata_pre_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!av_readdata_pre_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!av_readdata_pre_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!av_readdata_pre_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!av_readdata_pre_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!av_readdata_pre_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!av_readdata_pre_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!av_readdata_pre_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!av_readdata_pre_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!av_readdata_pre_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!av_readdata_pre_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!av_readdata_pre_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!av_readdata_pre_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!av_readdata_pre_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_1 (
	out_valid_reg,
	in_ready_hold,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_59,
	local_write,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	mem_116_0,
	mem_used_0,
	mem_59_0,
	mem_57_0,
	comb,
	mem_117_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	mem_100_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	in_data_reg_60,
	WideOr01,
	read,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	rp_valid,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
input 	in_ready_hold;
output 	mem_used_1;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
input 	local_write;
output 	write;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_116_0;
output 	mem_used_0;
output 	mem_59_0;
output 	mem_57_0;
input 	comb;
output 	mem_117_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	mem_100_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	in_data_reg_60;
input 	WideOr01;
output 	read;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_6;
input 	rp_valid;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;
input 	in_data_reg_100;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~1_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][116]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][59]~q ;
wire \mem~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem[1][117]~q ;
wire \mem~2_combout ;
wire \mem[1][69]~q ;
wire \mem~3_combout ;
wire \mem[1][68]~q ;
wire \mem~4_combout ;
wire \mem[1][67]~q ;
wire \mem~5_combout ;
wire \mem[1][66]~q ;
wire \mem~6_combout ;
wire \mem[1][65]~q ;
wire \mem~7_combout ;
wire \mem[1][92]~q ;
wire \mem~8_combout ;
wire \mem[1][93]~q ;
wire \mem~9_combout ;
wire \mem[1][94]~q ;
wire \mem~10_combout ;
wire \mem[1][95]~q ;
wire \mem~11_combout ;
wire \mem[1][96]~q ;
wire \mem~12_combout ;
wire \mem[1][97]~q ;
wire \mem~13_combout ;
wire \mem[1][98]~q ;
wire \mem~14_combout ;
wire \mem[1][99]~q ;
wire \mem~15_combout ;
wire \mem[1][100]~q ;
wire \mem~16_combout ;
wire \mem[1][101]~q ;
wire \mem~17_combout ;
wire \mem[1][102]~q ;
wire \mem~18_combout ;
wire \mem[1][103]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!in_ready_hold),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!local_write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \write~0 .shared_arith = "off";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][117] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_117_0),
	.prn(vcc));
defparam \mem[0][117] .is_wysiwyg = "true";
defparam \mem[0][117] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

dffeas \mem[0][100] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_100_0),
	.prn(vcc));
defparam \mem[0][100] .is_wysiwyg = "true";
defparam \mem[0][100] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!in_data_reg_59),
	.datab(!out_valid_reg),
	.datac(!write),
	.datad(!nxt_out_eop),
	.datae(!in_data_reg_60),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0001030300010303;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!\write~1_combout ),
	.datae(!read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5533055355330553;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][116]~q ),
	.datad(!in_data_reg_59),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_60),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!\write~1_combout ),
	.dataf(!read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3333FFFF1333FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][117] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][117]~q ),
	.prn(vcc));
defparam \mem[1][117] .is_wysiwyg = "true";
defparam \mem[1][117] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][117]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][100] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][100]~q ),
	.prn(vcc));
defparam \mem[1][100] .is_wysiwyg = "true";
defparam \mem[1][100] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][100]~q ),
	.datac(!in_data_reg_100),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_2 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_9,
	mem_9_0,
	av_readdata_pre_10,
	mem_10_0,
	av_readdata_pre_11,
	mem_11_0,
	av_readdata_pre_12,
	mem_12_0,
	av_readdata_pre_13,
	mem_13_0,
	av_readdata_pre_14,
	mem_14_0,
	av_readdata_pre_15,
	mem_15_0,
	av_readdata_pre_16,
	mem_16_0,
	av_readdata_pre_17,
	mem_17_0,
	av_readdata_pre_18,
	mem_18_0,
	av_readdata_pre_19,
	mem_19_0,
	av_readdata_pre_20,
	mem_20_0,
	av_readdata_pre_21,
	mem_21_0,
	av_readdata_pre_22,
	mem_22_0,
	av_readdata_pre_23,
	mem_23_0,
	av_readdata_pre_24,
	mem_24_0,
	av_readdata_pre_25,
	mem_25_0,
	av_readdata_pre_26,
	mem_26_0,
	av_readdata_pre_27,
	mem_27_0,
	av_readdata_pre_28,
	mem_28_0,
	av_readdata_pre_29,
	mem_29_0,
	av_readdata_pre_30,
	mem_30_0,
	av_readdata_pre_31,
	mem_31_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	always4;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	av_readdata_pre_8;
output 	mem_8_0;
input 	av_readdata_pre_9;
output 	mem_9_0;
input 	av_readdata_pre_10;
output 	mem_10_0;
input 	av_readdata_pre_11;
output 	mem_11_0;
input 	av_readdata_pre_12;
output 	mem_12_0;
input 	av_readdata_pre_13;
output 	mem_13_0;
input 	av_readdata_pre_14;
output 	mem_14_0;
input 	av_readdata_pre_15;
output 	mem_15_0;
input 	av_readdata_pre_16;
output 	mem_16_0;
input 	av_readdata_pre_17;
output 	mem_17_0;
input 	av_readdata_pre_18;
output 	mem_18_0;
input 	av_readdata_pre_19;
output 	mem_19_0;
input 	av_readdata_pre_20;
output 	mem_20_0;
input 	av_readdata_pre_21;
output 	mem_21_0;
input 	av_readdata_pre_22;
output 	mem_22_0;
input 	av_readdata_pre_23;
output 	mem_23_0;
input 	av_readdata_pre_24;
output 	mem_24_0;
input 	av_readdata_pre_25;
output 	mem_25_0;
input 	av_readdata_pre_26;
output 	mem_26_0;
input 	av_readdata_pre_27;
output 	mem_27_0;
input 	av_readdata_pre_28;
output 	mem_28_0;
input 	av_readdata_pre_29;
output 	mem_29_0;
input 	av_readdata_pre_30;
output 	mem_30_0;
input 	av_readdata_pre_31;
output 	mem_31_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!av_readdata_pre_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!av_readdata_pre_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!av_readdata_pre_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!av_readdata_pre_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!av_readdata_pre_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!av_readdata_pre_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!av_readdata_pre_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!av_readdata_pre_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!av_readdata_pre_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!av_readdata_pre_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!av_readdata_pre_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!av_readdata_pre_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!av_readdata_pre_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!av_readdata_pre_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!av_readdata_pre_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!av_readdata_pre_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!av_readdata_pre_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!av_readdata_pre_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!av_readdata_pre_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!av_readdata_pre_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!av_readdata_pre_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!av_readdata_pre_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_3 (
	in_ready_hold,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_59,
	local_write,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	mem_116_0,
	mem_used_0,
	mem_59_0,
	mem_57_0,
	comb,
	mem_117_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	mem_100_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	in_data_reg_60,
	WideOr01,
	read,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	rp_valid,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
input 	local_write;
output 	write;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_116_0;
output 	mem_used_0;
output 	mem_59_0;
output 	mem_57_0;
input 	comb;
output 	mem_117_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	mem_100_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	in_data_reg_60;
input 	WideOr01;
output 	read;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_6;
input 	rp_valid;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;
input 	in_data_reg_100;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~1_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][116]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][59]~q ;
wire \mem~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem[1][117]~q ;
wire \mem~2_combout ;
wire \mem[1][69]~q ;
wire \mem~3_combout ;
wire \mem[1][68]~q ;
wire \mem~4_combout ;
wire \mem[1][67]~q ;
wire \mem~5_combout ;
wire \mem[1][66]~q ;
wire \mem~6_combout ;
wire \mem[1][65]~q ;
wire \mem~7_combout ;
wire \mem[1][92]~q ;
wire \mem~8_combout ;
wire \mem[1][93]~q ;
wire \mem~9_combout ;
wire \mem[1][94]~q ;
wire \mem~10_combout ;
wire \mem[1][95]~q ;
wire \mem~11_combout ;
wire \mem[1][96]~q ;
wire \mem~12_combout ;
wire \mem[1][97]~q ;
wire \mem~13_combout ;
wire \mem[1][98]~q ;
wire \mem~14_combout ;
wire \mem[1][99]~q ;
wire \mem~15_combout ;
wire \mem[1][100]~q ;
wire \mem~16_combout ;
wire \mem[1][101]~q ;
wire \mem~17_combout ;
wire \mem[1][102]~q ;
wire \mem~18_combout ;
wire \mem[1][103]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!in_ready_hold),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!local_write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \write~0 .shared_arith = "off";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][117] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_117_0),
	.prn(vcc));
defparam \mem[0][117] .is_wysiwyg = "true";
defparam \mem[0][117] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

dffeas \mem[0][100] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_100_0),
	.prn(vcc));
defparam \mem[0][100] .is_wysiwyg = "true";
defparam \mem[0][100] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!in_data_reg_59),
	.datab(!out_valid_reg),
	.datac(!write),
	.datad(!nxt_out_eop),
	.datae(!in_data_reg_60),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0001030300010303;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!\write~1_combout ),
	.datae(!read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5533055355330553;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][116]~q ),
	.datad(!in_data_reg_59),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_60),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!\write~1_combout ),
	.dataf(!read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3333FFFF1333FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][117] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][117]~q ),
	.prn(vcc));
defparam \mem[1][117] .is_wysiwyg = "true";
defparam \mem[1][117] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][117]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][100] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][100]~q ),
	.prn(vcc));
defparam \mem[1][100] .is_wysiwyg = "true";
defparam \mem[1][100] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][100]~q ),
	.datac(!in_data_reg_100),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_4 (
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_9,
	mem_9_0,
	reset,
	WideOr0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	av_readdata_pre_0;
output 	always4;
output 	mem_0_0;
input 	av_readdata_pre_1;
output 	mem_1_0;
input 	av_readdata_pre_2;
output 	mem_2_0;
input 	av_readdata_pre_3;
output 	mem_3_0;
input 	av_readdata_pre_4;
output 	mem_4_0;
input 	av_readdata_pre_5;
output 	mem_5_0;
input 	av_readdata_pre_6;
output 	mem_6_0;
input 	av_readdata_pre_7;
output 	mem_7_0;
input 	av_readdata_pre_8;
output 	mem_8_0;
input 	av_readdata_pre_9;
output 	mem_9_0;
input 	reset;
input 	WideOr0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always4),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h4444444444444444;
defparam \always4~0 .shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!WideOr0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h0000777000007770;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h1F001F001F001F00;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!\mem_used[1]~q ),
	.datad(!\read~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h731F731F731F731F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!\read~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_5 (
	in_ready_hold,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_59,
	local_write,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	mem_116_0,
	mem_used_0,
	mem_59_0,
	mem_57_0,
	comb,
	mem_117_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	mem_100_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	in_data_reg_60,
	WideOr01,
	read,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	rp_valid,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	out_valid_reg;
output 	mem_used_1;
input 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
input 	local_write;
output 	write;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_116_0;
output 	mem_used_0;
output 	mem_59_0;
output 	mem_57_0;
input 	comb;
output 	mem_117_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	mem_100_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	in_data_reg_60;
input 	WideOr01;
output 	read;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_6;
input 	rp_valid;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;
input 	in_data_reg_100;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~1_combout ;
wire \mem_used[1]~0_combout ;
wire \mem[1][116]~q ;
wire \mem~20_combout ;
wire \always0~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][59]~q ;
wire \mem~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem[1][117]~q ;
wire \mem~2_combout ;
wire \mem[1][69]~q ;
wire \mem~3_combout ;
wire \mem[1][68]~q ;
wire \mem~4_combout ;
wire \mem[1][67]~q ;
wire \mem~5_combout ;
wire \mem[1][66]~q ;
wire \mem~6_combout ;
wire \mem[1][65]~q ;
wire \mem~7_combout ;
wire \mem[1][92]~q ;
wire \mem~8_combout ;
wire \mem[1][93]~q ;
wire \mem~9_combout ;
wire \mem[1][94]~q ;
wire \mem~10_combout ;
wire \mem[1][95]~q ;
wire \mem~11_combout ;
wire \mem[1][96]~q ;
wire \mem~12_combout ;
wire \mem[1][97]~q ;
wire \mem~13_combout ;
wire \mem[1][98]~q ;
wire \mem~14_combout ;
wire \mem[1][99]~q ;
wire \mem~15_combout ;
wire \mem[1][100]~q ;
wire \mem~16_combout ;
wire \mem[1][101]~q ;
wire \mem~17_combout ;
wire \mem[1][102]~q ;
wire \mem~18_combout ;
wire \mem[1][103]~q ;
wire \mem~19_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!in_ready_hold),
	.datab(!mem_used_1),
	.datac(!WideOr0),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(!local_write),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hC0C0C4C0C4C0C0C0;
defparam \write~0 .shared_arith = "off";

dffeas \mem[0][116] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_116_0),
	.prn(vcc));
defparam \mem[0][116] .is_wysiwyg = "true";
defparam \mem[0][116] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_59_0),
	.prn(vcc));
defparam \mem[0][59] .is_wysiwyg = "true";
defparam \mem[0][59] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem[0][117] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_117_0),
	.prn(vcc));
defparam \mem[0][117] .is_wysiwyg = "true";
defparam \mem[0][117] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

dffeas \mem[0][100] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_100_0),
	.prn(vcc));
defparam \mem[0][100] .is_wysiwyg = "true";
defparam \mem[0][100] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!comb),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h1111111111111111;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!in_data_reg_59),
	.datab(!out_valid_reg),
	.datac(!write),
	.datad(!nxt_out_eop),
	.datae(!in_data_reg_60),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0001030300010303;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!\write~1_combout ),
	.datae(!read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5533055355330553;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][116] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][116]~q ),
	.prn(vcc));
defparam \mem[1][116] .is_wysiwyg = "true";
defparam \mem[1][116] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!WideOr0),
	.datab(!out_valid_reg),
	.datac(!\mem[1][116]~q ),
	.datad(!in_data_reg_59),
	.datae(!mem_used_1),
	.dataf(!nxt_out_eop),
	.datag(!in_data_reg_60),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "on";
defparam \mem~20 .lut_mask = 64'h02020F0F02330F0F;
defparam \mem~20 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!rp_valid),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAAEAAAEAAAEAAAEA;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!rp_valid),
	.datad(!last_packet_beat),
	.datae(!\write~1_combout ),
	.dataf(!read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3333FFFF1333FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][59] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][59]~q ),
	.prn(vcc));
defparam \mem[1][59] .is_wysiwyg = "true";
defparam \mem[1][59] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_59),
	.datac(!\mem[1][59]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][117] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][117]~q ),
	.prn(vcc));
defparam \mem[1][117] .is_wysiwyg = "true";
defparam \mem[1][117] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][117]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h2727272727272727;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h0257025702570257;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][100] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][100]~q ),
	.prn(vcc));
defparam \mem[1][100] .is_wysiwyg = "true";
defparam \mem[1][100] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][100]~q ),
	.datac(!in_data_reg_100),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~19 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_6 (
	h2f_lw_RREADY_0,
	in_ready_hold,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	mem_11_0,
	av_readdata_pre_30,
	mem_10_0,
	reset,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_RREADY_0;
input 	in_ready_hold;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
output 	mem_11_0;
input 	av_readdata_pre_30;
output 	mem_10_0;
input 	reset;
output 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][30]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][10]~q ;
wire \mem~1_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!empty1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4444444444444444;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!in_ready_hold),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_7 (
	in_ready_hold,
	mem_used_1,
	in_data_reg_60,
	wait_latency_counter_1,
	wait_latency_counter_0,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_117_0,
	mem_57_0,
	mem_used_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	mem_100_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	read,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
output 	mem_used_1;
input 	in_data_reg_60;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_117_0;
output 	mem_57_0;
output 	mem_used_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	mem_100_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	read;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;
input 	in_data_reg_100;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~0_combout ;
wire \mem[1][117]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][69]~q ;
wire \mem~2_combout ;
wire \mem[1][68]~q ;
wire \mem~3_combout ;
wire \mem[1][67]~q ;
wire \mem~4_combout ;
wire \mem[1][66]~q ;
wire \mem~5_combout ;
wire \mem[1][65]~q ;
wire \mem~6_combout ;
wire \mem[1][92]~q ;
wire \mem~7_combout ;
wire \mem[1][93]~q ;
wire \mem~8_combout ;
wire \mem[1][94]~q ;
wire \mem~9_combout ;
wire \mem[1][95]~q ;
wire \mem~10_combout ;
wire \mem[1][96]~q ;
wire \mem~11_combout ;
wire \mem[1][97]~q ;
wire \mem~12_combout ;
wire \mem[1][98]~q ;
wire \mem~13_combout ;
wire \mem[1][99]~q ;
wire \mem~14_combout ;
wire \mem[1][100]~q ;
wire \mem~15_combout ;
wire \mem[1][101]~q ;
wire \mem~16_combout ;
wire \mem[1][102]~q ;
wire \mem~17_combout ;
wire \mem[1][103]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][117] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_117_0),
	.prn(vcc));
defparam \mem[0][117] .is_wysiwyg = "true";
defparam \mem[0][117] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

dffeas \mem[0][100] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_100_0),
	.prn(vcc));
defparam \mem[0][100] .is_wysiwyg = "true";
defparam \mem[0][100] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!in_ready_hold),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0002000200020002;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5545331355453313;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][117] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][117]~q ),
	.prn(vcc));
defparam \mem[1][117] .is_wysiwyg = "true";
defparam \mem[1][117] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][117]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!last_packet_beat),
	.datac(!read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAEAEAEAEAEAEAEAE;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3313FFFF3313FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][100] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][100]~q ),
	.prn(vcc));
defparam \mem[1][100] .is_wysiwyg = "true";
defparam \mem[1][100] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][100]~q ),
	.datac(!in_data_reg_100),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_8 (
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	mem_0_0,
	av_readdata_pre_0,
	mem_1_0,
	av_readdata_pre_1,
	mem_2_0,
	av_readdata_pre_2,
	mem_3_0,
	av_readdata_pre_3,
	mem_4_0,
	av_readdata_pre_4,
	mem_5_0,
	av_readdata_pre_5,
	mem_6_0,
	av_readdata_pre_6,
	mem_7_0,
	av_readdata_pre_7,
	mem_8_0,
	av_readdata_pre_8,
	av_readdata_pre_9,
	mem_9_0,
	mem_10_0,
	av_readdata_pre_10,
	mem_11_0,
	av_readdata_pre_11,
	mem_12_0,
	av_readdata_pre_12,
	mem_13_0,
	av_readdata_pre_13,
	mem_14_0,
	av_readdata_pre_14,
	mem_15_0,
	av_readdata_pre_15,
	mem_16_0,
	av_readdata_pre_16,
	mem_17_0,
	av_readdata_pre_17,
	mem_18_0,
	av_readdata_pre_18,
	mem_19_0,
	av_readdata_pre_19,
	mem_20_0,
	av_readdata_pre_20,
	mem_21_0,
	av_readdata_pre_21,
	mem_22_0,
	av_readdata_pre_22,
	mem_23_0,
	av_readdata_pre_23,
	mem_24_0,
	av_readdata_pre_24,
	mem_25_0,
	av_readdata_pre_25,
	mem_26_0,
	av_readdata_pre_26,
	mem_27_0,
	av_readdata_pre_27,
	mem_28_0,
	av_readdata_pre_28,
	mem_29_0,
	av_readdata_pre_29,
	mem_30_0,
	av_readdata_pre_30,
	mem_31_0,
	av_readdata_pre_31,
	reset,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
output 	mem_0_0;
input 	av_readdata_pre_0;
output 	mem_1_0;
input 	av_readdata_pre_1;
output 	mem_2_0;
input 	av_readdata_pre_2;
output 	mem_3_0;
input 	av_readdata_pre_3;
output 	mem_4_0;
input 	av_readdata_pre_4;
output 	mem_5_0;
input 	av_readdata_pre_5;
output 	mem_6_0;
input 	av_readdata_pre_6;
output 	mem_7_0;
input 	av_readdata_pre_7;
output 	mem_8_0;
input 	av_readdata_pre_8;
input 	av_readdata_pre_9;
output 	mem_9_0;
output 	mem_10_0;
input 	av_readdata_pre_10;
output 	mem_11_0;
input 	av_readdata_pre_11;
output 	mem_12_0;
input 	av_readdata_pre_12;
output 	mem_13_0;
input 	av_readdata_pre_13;
output 	mem_14_0;
input 	av_readdata_pre_14;
output 	mem_15_0;
input 	av_readdata_pre_15;
output 	mem_16_0;
input 	av_readdata_pre_16;
output 	mem_17_0;
input 	av_readdata_pre_17;
output 	mem_18_0;
input 	av_readdata_pre_18;
output 	mem_19_0;
input 	av_readdata_pre_19;
output 	mem_20_0;
input 	av_readdata_pre_20;
output 	mem_21_0;
input 	av_readdata_pre_21;
output 	mem_22_0;
input 	av_readdata_pre_22;
output 	mem_23_0;
input 	av_readdata_pre_23;
output 	mem_24_0;
input 	av_readdata_pre_24;
output 	mem_25_0;
input 	av_readdata_pre_25;
output 	mem_26_0;
input 	av_readdata_pre_26;
output 	mem_27_0;
input 	av_readdata_pre_27;
output 	mem_28_0;
input 	av_readdata_pre_28;
output 	mem_29_0;
input 	av_readdata_pre_29;
output 	mem_30_0;
input 	av_readdata_pre_30;
output 	mem_31_0;
input 	av_readdata_pre_31;
input 	reset;
output 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;
wire \mem[1][10]~q ;
wire \mem~10_combout ;
wire \mem[1][11]~q ;
wire \mem~11_combout ;
wire \mem[1][12]~q ;
wire \mem~12_combout ;
wire \mem[1][13]~q ;
wire \mem~13_combout ;
wire \mem[1][14]~q ;
wire \mem~14_combout ;
wire \mem[1][15]~q ;
wire \mem~15_combout ;
wire \mem[1][16]~q ;
wire \mem~16_combout ;
wire \mem[1][17]~q ;
wire \mem~17_combout ;
wire \mem[1][18]~q ;
wire \mem~18_combout ;
wire \mem[1][19]~q ;
wire \mem~19_combout ;
wire \mem[1][20]~q ;
wire \mem~20_combout ;
wire \mem[1][21]~q ;
wire \mem~21_combout ;
wire \mem[1][22]~q ;
wire \mem~22_combout ;
wire \mem[1][23]~q ;
wire \mem~23_combout ;
wire \mem[1][24]~q ;
wire \mem~24_combout ;
wire \mem[1][25]~q ;
wire \mem~25_combout ;
wire \mem[1][26]~q ;
wire \mem~26_combout ;
wire \mem[1][27]~q ;
wire \mem~27_combout ;
wire \mem[1][28]~q ;
wire \mem~28_combout ;
wire \mem[1][29]~q ;
wire \mem~29_combout ;
wire \mem[1][30]~q ;
wire \mem~30_combout ;
wire \mem[1][31]~q ;
wire \mem~31_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

dffeas \mem[0][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_10_0),
	.prn(vcc));
defparam \mem[0][10] .is_wysiwyg = "true";
defparam \mem[0][10] .power_up = "low";

dffeas \mem[0][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_11_0),
	.prn(vcc));
defparam \mem[0][11] .is_wysiwyg = "true";
defparam \mem[0][11] .power_up = "low";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_12_0),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[0][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_13_0),
	.prn(vcc));
defparam \mem[0][13] .is_wysiwyg = "true";
defparam \mem[0][13] .power_up = "low";

dffeas \mem[0][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_14_0),
	.prn(vcc));
defparam \mem[0][14] .is_wysiwyg = "true";
defparam \mem[0][14] .power_up = "low";

dffeas \mem[0][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_15_0),
	.prn(vcc));
defparam \mem[0][15] .is_wysiwyg = "true";
defparam \mem[0][15] .power_up = "low";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_16_0),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[0][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_17_0),
	.prn(vcc));
defparam \mem[0][17] .is_wysiwyg = "true";
defparam \mem[0][17] .power_up = "low";

dffeas \mem[0][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_18_0),
	.prn(vcc));
defparam \mem[0][18] .is_wysiwyg = "true";
defparam \mem[0][18] .power_up = "low";

dffeas \mem[0][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_19_0),
	.prn(vcc));
defparam \mem[0][19] .is_wysiwyg = "true";
defparam \mem[0][19] .power_up = "low";

dffeas \mem[0][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_20_0),
	.prn(vcc));
defparam \mem[0][20] .is_wysiwyg = "true";
defparam \mem[0][20] .power_up = "low";

dffeas \mem[0][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_21_0),
	.prn(vcc));
defparam \mem[0][21] .is_wysiwyg = "true";
defparam \mem[0][21] .power_up = "low";

dffeas \mem[0][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_22_0),
	.prn(vcc));
defparam \mem[0][22] .is_wysiwyg = "true";
defparam \mem[0][22] .power_up = "low";

dffeas \mem[0][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_23_0),
	.prn(vcc));
defparam \mem[0][23] .is_wysiwyg = "true";
defparam \mem[0][23] .power_up = "low";

dffeas \mem[0][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_24_0),
	.prn(vcc));
defparam \mem[0][24] .is_wysiwyg = "true";
defparam \mem[0][24] .power_up = "low";

dffeas \mem[0][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_25_0),
	.prn(vcc));
defparam \mem[0][25] .is_wysiwyg = "true";
defparam \mem[0][25] .power_up = "low";

dffeas \mem[0][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_26_0),
	.prn(vcc));
defparam \mem[0][26] .is_wysiwyg = "true";
defparam \mem[0][26] .power_up = "low";

dffeas \mem[0][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_27_0),
	.prn(vcc));
defparam \mem[0][27] .is_wysiwyg = "true";
defparam \mem[0][27] .power_up = "low";

dffeas \mem[0][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_28_0),
	.prn(vcc));
defparam \mem[0][28] .is_wysiwyg = "true";
defparam \mem[0][28] .power_up = "low";

dffeas \mem[0][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_29_0),
	.prn(vcc));
defparam \mem[0][29] .is_wysiwyg = "true";
defparam \mem[0][29] .power_up = "low";

dffeas \mem[0][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_30_0),
	.prn(vcc));
defparam \mem[0][30] .is_wysiwyg = "true";
defparam \mem[0][30] .power_up = "low";

dffeas \mem[0][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_31_0),
	.prn(vcc));
defparam \mem[0][31] .is_wysiwyg = "true";
defparam \mem[0][31] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!empty1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4444444444444444;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][10] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][10]~q ),
	.prn(vcc));
defparam \mem[1][10] .is_wysiwyg = "true";
defparam \mem[1][10] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!av_readdata_pre_10),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h4747474747474747;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][11] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][11]~q ),
	.prn(vcc));
defparam \mem[1][11] .is_wysiwyg = "true";
defparam \mem[1][11] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!av_readdata_pre_11),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h4747474747474747;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!av_readdata_pre_12),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h4747474747474747;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][13] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][13]~q ),
	.prn(vcc));
defparam \mem[1][13] .is_wysiwyg = "true";
defparam \mem[1][13] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!av_readdata_pre_13),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h4747474747474747;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][14] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][14]~q ),
	.prn(vcc));
defparam \mem[1][14] .is_wysiwyg = "true";
defparam \mem[1][14] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!av_readdata_pre_14),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h4747474747474747;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][15] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][15]~q ),
	.prn(vcc));
defparam \mem[1][15] .is_wysiwyg = "true";
defparam \mem[1][15] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!av_readdata_pre_15),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h4747474747474747;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!av_readdata_pre_16),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h4747474747474747;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][17] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][17]~q ),
	.prn(vcc));
defparam \mem[1][17] .is_wysiwyg = "true";
defparam \mem[1][17] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!av_readdata_pre_17),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h4747474747474747;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][18] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][18]~q ),
	.prn(vcc));
defparam \mem[1][18] .is_wysiwyg = "true";
defparam \mem[1][18] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!av_readdata_pre_18),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h4747474747474747;
defparam \mem~18 .shared_arith = "off";

dffeas \mem[1][19] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][19]~q ),
	.prn(vcc));
defparam \mem[1][19] .is_wysiwyg = "true";
defparam \mem[1][19] .power_up = "low";

cyclonev_lcell_comb \mem~19 (
	.dataa(!av_readdata_pre_19),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~19 .extended_lut = "off";
defparam \mem~19 .lut_mask = 64'h4747474747474747;
defparam \mem~19 .shared_arith = "off";

dffeas \mem[1][20] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][20]~q ),
	.prn(vcc));
defparam \mem[1][20] .is_wysiwyg = "true";
defparam \mem[1][20] .power_up = "low";

cyclonev_lcell_comb \mem~20 (
	.dataa(!av_readdata_pre_20),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~20 .extended_lut = "off";
defparam \mem~20 .lut_mask = 64'h4747474747474747;
defparam \mem~20 .shared_arith = "off";

dffeas \mem[1][21] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][21]~q ),
	.prn(vcc));
defparam \mem[1][21] .is_wysiwyg = "true";
defparam \mem[1][21] .power_up = "low";

cyclonev_lcell_comb \mem~21 (
	.dataa(!av_readdata_pre_21),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~21 .extended_lut = "off";
defparam \mem~21 .lut_mask = 64'h4747474747474747;
defparam \mem~21 .shared_arith = "off";

dffeas \mem[1][22] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][22]~q ),
	.prn(vcc));
defparam \mem[1][22] .is_wysiwyg = "true";
defparam \mem[1][22] .power_up = "low";

cyclonev_lcell_comb \mem~22 (
	.dataa(!av_readdata_pre_22),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~22 .extended_lut = "off";
defparam \mem~22 .lut_mask = 64'h4747474747474747;
defparam \mem~22 .shared_arith = "off";

dffeas \mem[1][23] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][23]~q ),
	.prn(vcc));
defparam \mem[1][23] .is_wysiwyg = "true";
defparam \mem[1][23] .power_up = "low";

cyclonev_lcell_comb \mem~23 (
	.dataa(!av_readdata_pre_23),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~23 .extended_lut = "off";
defparam \mem~23 .lut_mask = 64'h4747474747474747;
defparam \mem~23 .shared_arith = "off";

dffeas \mem[1][24] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][24]~q ),
	.prn(vcc));
defparam \mem[1][24] .is_wysiwyg = "true";
defparam \mem[1][24] .power_up = "low";

cyclonev_lcell_comb \mem~24 (
	.dataa(!av_readdata_pre_24),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~24 .extended_lut = "off";
defparam \mem~24 .lut_mask = 64'h4747474747474747;
defparam \mem~24 .shared_arith = "off";

dffeas \mem[1][25] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][25]~q ),
	.prn(vcc));
defparam \mem[1][25] .is_wysiwyg = "true";
defparam \mem[1][25] .power_up = "low";

cyclonev_lcell_comb \mem~25 (
	.dataa(!av_readdata_pre_25),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~25 .extended_lut = "off";
defparam \mem~25 .lut_mask = 64'h4747474747474747;
defparam \mem~25 .shared_arith = "off";

dffeas \mem[1][26] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][26]~q ),
	.prn(vcc));
defparam \mem[1][26] .is_wysiwyg = "true";
defparam \mem[1][26] .power_up = "low";

cyclonev_lcell_comb \mem~26 (
	.dataa(!av_readdata_pre_26),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~26 .extended_lut = "off";
defparam \mem~26 .lut_mask = 64'h4747474747474747;
defparam \mem~26 .shared_arith = "off";

dffeas \mem[1][27] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][27]~q ),
	.prn(vcc));
defparam \mem[1][27] .is_wysiwyg = "true";
defparam \mem[1][27] .power_up = "low";

cyclonev_lcell_comb \mem~27 (
	.dataa(!av_readdata_pre_27),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~27 .extended_lut = "off";
defparam \mem~27 .lut_mask = 64'h4747474747474747;
defparam \mem~27 .shared_arith = "off";

dffeas \mem[1][28] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][28]~q ),
	.prn(vcc));
defparam \mem[1][28] .is_wysiwyg = "true";
defparam \mem[1][28] .power_up = "low";

cyclonev_lcell_comb \mem~28 (
	.dataa(!av_readdata_pre_28),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~28 .extended_lut = "off";
defparam \mem~28 .lut_mask = 64'h4747474747474747;
defparam \mem~28 .shared_arith = "off";

dffeas \mem[1][29] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][29]~q ),
	.prn(vcc));
defparam \mem[1][29] .is_wysiwyg = "true";
defparam \mem[1][29] .power_up = "low";

cyclonev_lcell_comb \mem~29 (
	.dataa(!av_readdata_pre_29),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~29 .extended_lut = "off";
defparam \mem~29 .lut_mask = 64'h4747474747474747;
defparam \mem~29 .shared_arith = "off";

dffeas \mem[1][30] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][30]~q ),
	.prn(vcc));
defparam \mem[1][30] .is_wysiwyg = "true";
defparam \mem[1][30] .power_up = "low";

cyclonev_lcell_comb \mem~30 (
	.dataa(!av_readdata_pre_30),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~30 .extended_lut = "off";
defparam \mem~30 .lut_mask = 64'h4747474747474747;
defparam \mem~30 .shared_arith = "off";

dffeas \mem[1][31] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][31]~q ),
	.prn(vcc));
defparam \mem[1][31] .is_wysiwyg = "true";
defparam \mem[1][31] .power_up = "low";

cyclonev_lcell_comb \mem~31 (
	.dataa(!av_readdata_pre_31),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~31 .extended_lut = "off";
defparam \mem~31 .lut_mask = 64'h4747474747474747;
defparam \mem~31 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_9 (
	in_ready_hold,
	mem_used_1,
	in_data_reg_60,
	wait_latency_counter_1,
	wait_latency_counter_0,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_117_0,
	mem_57_0,
	mem_used_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	mem_100_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	read,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
output 	mem_used_1;
input 	in_data_reg_60;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_117_0;
output 	mem_57_0;
output 	mem_used_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	mem_100_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	read;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;
input 	in_data_reg_100;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~0_combout ;
wire \mem[1][117]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][69]~q ;
wire \mem~2_combout ;
wire \mem[1][68]~q ;
wire \mem~3_combout ;
wire \mem[1][67]~q ;
wire \mem~4_combout ;
wire \mem[1][66]~q ;
wire \mem~5_combout ;
wire \mem[1][65]~q ;
wire \mem~6_combout ;
wire \mem[1][92]~q ;
wire \mem~7_combout ;
wire \mem[1][93]~q ;
wire \mem~8_combout ;
wire \mem[1][94]~q ;
wire \mem~9_combout ;
wire \mem[1][95]~q ;
wire \mem~10_combout ;
wire \mem[1][96]~q ;
wire \mem~11_combout ;
wire \mem[1][97]~q ;
wire \mem~12_combout ;
wire \mem[1][98]~q ;
wire \mem~13_combout ;
wire \mem[1][99]~q ;
wire \mem~14_combout ;
wire \mem[1][100]~q ;
wire \mem~15_combout ;
wire \mem[1][101]~q ;
wire \mem~16_combout ;
wire \mem[1][102]~q ;
wire \mem~17_combout ;
wire \mem[1][103]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][117] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_117_0),
	.prn(vcc));
defparam \mem[0][117] .is_wysiwyg = "true";
defparam \mem[0][117] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

dffeas \mem[0][100] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_100_0),
	.prn(vcc));
defparam \mem[0][100] .is_wysiwyg = "true";
defparam \mem[0][100] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!in_ready_hold),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0002000200020002;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5545331355453313;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][117] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][117]~q ),
	.prn(vcc));
defparam \mem[1][117] .is_wysiwyg = "true";
defparam \mem[1][117] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][117]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!last_packet_beat),
	.datac(!read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAEAEAEAEAEAEAEAE;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3313FFFF3313FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][100] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][100]~q ),
	.prn(vcc));
defparam \mem[1][100] .is_wysiwyg = "true";
defparam \mem[1][100] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][100]~q ),
	.datac(!in_data_reg_100),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_10 (
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	empty1,
	mem_0_0,
	av_readdata_pre_0,
	mem_1_0,
	av_readdata_pre_1,
	mem_2_0,
	av_readdata_pre_2,
	mem_3_0,
	av_readdata_pre_3,
	mem_4_0,
	av_readdata_pre_4,
	mem_5_0,
	av_readdata_pre_5,
	mem_6_0,
	av_readdata_pre_6,
	mem_7_0,
	av_readdata_pre_7,
	mem_8_0,
	av_readdata_pre_8,
	mem_9_0,
	av_readdata_pre_9,
	reset,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
output 	mem_used_0;
output 	empty1;
output 	mem_0_0;
input 	av_readdata_pre_0;
output 	mem_1_0;
input 	av_readdata_pre_1;
output 	mem_2_0;
input 	av_readdata_pre_2;
output 	mem_3_0;
input 	av_readdata_pre_3;
output 	mem_4_0;
input 	av_readdata_pre_4;
output 	mem_5_0;
input 	av_readdata_pre_5;
output 	mem_6_0;
input 	av_readdata_pre_6;
output 	mem_7_0;
input 	av_readdata_pre_7;
output 	mem_8_0;
input 	av_readdata_pre_8;
output 	mem_9_0;
input 	av_readdata_pre_9;
input 	reset;
output 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~1_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~0_combout ;
wire \mem[1][0]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][1]~q ;
wire \mem~1_combout ;
wire \mem[1][2]~q ;
wire \mem~2_combout ;
wire \mem[1][3]~q ;
wire \mem~3_combout ;
wire \mem[1][4]~q ;
wire \mem~4_combout ;
wire \mem[1][5]~q ;
wire \mem~5_combout ;
wire \mem[1][6]~q ;
wire \mem~6_combout ;
wire \mem[1][7]~q ;
wire \mem~7_combout ;
wire \mem[1][8]~q ;
wire \mem~8_combout ;
wire \mem[1][9]~q ;
wire \mem~9_combout ;


dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb empty(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(empty1),
	.sumout(),
	.cout(),
	.shareout());
defparam empty.extended_lut = "off";
defparam empty.lut_mask = 64'h8888888888888888;
defparam empty.shared_arith = "off";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_0_0),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_1_0),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_2_0),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[0][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_3_0),
	.prn(vcc));
defparam \mem[0][3] .is_wysiwyg = "true";
defparam \mem[0][3] .power_up = "low";

dffeas \mem[0][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_4_0),
	.prn(vcc));
defparam \mem[0][4] .is_wysiwyg = "true";
defparam \mem[0][4] .power_up = "low";

dffeas \mem[0][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_5_0),
	.prn(vcc));
defparam \mem[0][5] .is_wysiwyg = "true";
defparam \mem[0][5] .power_up = "low";

dffeas \mem[0][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_6_0),
	.prn(vcc));
defparam \mem[0][6] .is_wysiwyg = "true";
defparam \mem[0][6] .power_up = "low";

dffeas \mem[0][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_7_0),
	.prn(vcc));
defparam \mem[0][7] .is_wysiwyg = "true";
defparam \mem[0][7] .power_up = "low";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_8_0),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

dffeas \mem[0][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_9_0),
	.prn(vcc));
defparam \mem[0][9] .is_wysiwyg = "true";
defparam \mem[0][9] .power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!empty1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'h4444444444444444;
defparam \read~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'h02EA02EA02EA02EA;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_0),
	.datad(!\mem_used[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~0 .extended_lut = "off";
defparam \mem_used[0]~0 .lut_mask = 64'h2B1F2B1F2B1F2B1F;
defparam \mem_used[0]~0 .shared_arith = "off";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!av_readdata_pre_0),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h4747474747474747;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!h2f_lw_RREADY_0),
	.datab(!mem_used_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!av_readdata_pre_1),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h4747474747474747;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!av_readdata_pre_2),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h4747474747474747;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][3] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][3]~q ),
	.prn(vcc));
defparam \mem[1][3] .is_wysiwyg = "true";
defparam \mem[1][3] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!av_readdata_pre_3),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h4747474747474747;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][4] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][4]~q ),
	.prn(vcc));
defparam \mem[1][4] .is_wysiwyg = "true";
defparam \mem[1][4] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!av_readdata_pre_4),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h4747474747474747;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][5] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][5]~q ),
	.prn(vcc));
defparam \mem[1][5] .is_wysiwyg = "true";
defparam \mem[1][5] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!av_readdata_pre_5),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h4747474747474747;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][6] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][6]~q ),
	.prn(vcc));
defparam \mem[1][6] .is_wysiwyg = "true";
defparam \mem[1][6] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!av_readdata_pre_6),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h4747474747474747;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][7] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][7]~q ),
	.prn(vcc));
defparam \mem[1][7] .is_wysiwyg = "true";
defparam \mem[1][7] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!av_readdata_pre_7),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h4747474747474747;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!av_readdata_pre_8),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h4747474747474747;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][9] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][9]~q ),
	.prn(vcc));
defparam \mem[1][9] .is_wysiwyg = "true";
defparam \mem[1][9] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!av_readdata_pre_9),
	.datab(!\mem_used[1]~q ),
	.datac(!\mem[1][9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h4747474747474747;
defparam \mem~9 .shared_arith = "off";

endmodule

module terminal_qsys_altera_avalon_sc_fifo_11 (
	mem_used_1,
	in_data_reg_60,
	in_ready_hold,
	wait_latency_counter_1,
	wait_latency_counter_0,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	mem_117_0,
	mem_57_0,
	mem_used_0,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	mem_92_0,
	mem_93_0,
	mem_94_0,
	mem_95_0,
	mem_96_0,
	mem_97_0,
	mem_98_0,
	mem_99_0,
	mem_100_0,
	mem_101_0,
	mem_102_0,
	mem_103_0,
	reset,
	nxt_out_eop,
	last_packet_beat,
	read,
	write,
	write1,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	clk)/* synthesis synthesis_greybox=0 */;
output 	mem_used_1;
input 	in_data_reg_60;
input 	in_ready_hold;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	out_valid_reg;
input 	stateST_UNCOMP_WR_SUBBURST;
output 	mem_117_0;
output 	mem_57_0;
output 	mem_used_0;
output 	mem_69_0;
output 	mem_68_0;
output 	mem_67_0;
output 	mem_66_0;
output 	mem_65_0;
output 	mem_92_0;
output 	mem_93_0;
output 	mem_94_0;
output 	mem_95_0;
output 	mem_96_0;
output 	mem_97_0;
output 	mem_98_0;
output 	mem_99_0;
output 	mem_100_0;
output 	mem_101_0;
output 	mem_102_0;
output 	mem_103_0;
input 	reset;
input 	nxt_out_eop;
input 	last_packet_beat;
input 	read;
output 	write;
output 	write1;
input 	out_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_5;
input 	out_uncomp_byte_cnt_reg_4;
input 	out_uncomp_byte_cnt_reg_3;
input 	out_uncomp_byte_cnt_reg_2;
input 	out_uncomp_byte_cnt_reg_6;
input 	in_data_reg_92;
input 	in_data_reg_93;
input 	in_data_reg_94;
input 	in_data_reg_95;
input 	in_data_reg_96;
input 	in_data_reg_97;
input 	in_data_reg_98;
input 	in_data_reg_99;
input 	in_data_reg_100;
input 	in_data_reg_101;
input 	in_data_reg_102;
input 	in_data_reg_103;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[1]~0_combout ;
wire \mem[1][117]~q ;
wire \mem~0_combout ;
wire \always0~0_combout ;
wire \mem[1][60]~q ;
wire \mem~1_combout ;
wire \mem_used[0]~1_combout ;
wire \mem[1][69]~q ;
wire \mem~2_combout ;
wire \mem[1][68]~q ;
wire \mem~3_combout ;
wire \mem[1][67]~q ;
wire \mem~4_combout ;
wire \mem[1][66]~q ;
wire \mem~5_combout ;
wire \mem[1][65]~q ;
wire \mem~6_combout ;
wire \mem[1][92]~q ;
wire \mem~7_combout ;
wire \mem[1][93]~q ;
wire \mem~8_combout ;
wire \mem[1][94]~q ;
wire \mem~9_combout ;
wire \mem[1][95]~q ;
wire \mem~10_combout ;
wire \mem[1][96]~q ;
wire \mem~11_combout ;
wire \mem[1][97]~q ;
wire \mem~12_combout ;
wire \mem[1][98]~q ;
wire \mem~13_combout ;
wire \mem[1][99]~q ;
wire \mem~14_combout ;
wire \mem[1][100]~q ;
wire \mem~15_combout ;
wire \mem[1][101]~q ;
wire \mem~16_combout ;
wire \mem[1][102]~q ;
wire \mem~17_combout ;
wire \mem[1][103]~q ;
wire \mem~18_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][117] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_117_0),
	.prn(vcc));
defparam \mem[0][117] .is_wysiwyg = "true";
defparam \mem[0][117] .power_up = "low";

dffeas \mem[0][57] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_57_0),
	.prn(vcc));
defparam \mem[0][57] .is_wysiwyg = "true";
defparam \mem[0][57] .power_up = "low";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_0),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

dffeas \mem[0][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_69_0),
	.prn(vcc));
defparam \mem[0][69] .is_wysiwyg = "true";
defparam \mem[0][69] .power_up = "low";

dffeas \mem[0][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_68_0),
	.prn(vcc));
defparam \mem[0][68] .is_wysiwyg = "true";
defparam \mem[0][68] .power_up = "low";

dffeas \mem[0][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_67_0),
	.prn(vcc));
defparam \mem[0][67] .is_wysiwyg = "true";
defparam \mem[0][67] .power_up = "low";

dffeas \mem[0][66] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_66_0),
	.prn(vcc));
defparam \mem[0][66] .is_wysiwyg = "true";
defparam \mem[0][66] .power_up = "low";

dffeas \mem[0][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_65_0),
	.prn(vcc));
defparam \mem[0][65] .is_wysiwyg = "true";
defparam \mem[0][65] .power_up = "low";

dffeas \mem[0][92] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_92_0),
	.prn(vcc));
defparam \mem[0][92] .is_wysiwyg = "true";
defparam \mem[0][92] .power_up = "low";

dffeas \mem[0][93] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_93_0),
	.prn(vcc));
defparam \mem[0][93] .is_wysiwyg = "true";
defparam \mem[0][93] .power_up = "low";

dffeas \mem[0][94] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_94_0),
	.prn(vcc));
defparam \mem[0][94] .is_wysiwyg = "true";
defparam \mem[0][94] .power_up = "low";

dffeas \mem[0][95] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_95_0),
	.prn(vcc));
defparam \mem[0][95] .is_wysiwyg = "true";
defparam \mem[0][95] .power_up = "low";

dffeas \mem[0][96] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_96_0),
	.prn(vcc));
defparam \mem[0][96] .is_wysiwyg = "true";
defparam \mem[0][96] .power_up = "low";

dffeas \mem[0][97] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_97_0),
	.prn(vcc));
defparam \mem[0][97] .is_wysiwyg = "true";
defparam \mem[0][97] .power_up = "low";

dffeas \mem[0][98] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_98_0),
	.prn(vcc));
defparam \mem[0][98] .is_wysiwyg = "true";
defparam \mem[0][98] .power_up = "low";

dffeas \mem[0][99] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_99_0),
	.prn(vcc));
defparam \mem[0][99] .is_wysiwyg = "true";
defparam \mem[0][99] .power_up = "low";

dffeas \mem[0][100] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_100_0),
	.prn(vcc));
defparam \mem[0][100] .is_wysiwyg = "true";
defparam \mem[0][100] .power_up = "low";

dffeas \mem[0][101] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_101_0),
	.prn(vcc));
defparam \mem[0][101] .is_wysiwyg = "true";
defparam \mem[0][101] .power_up = "low";

dffeas \mem[0][102] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_102_0),
	.prn(vcc));
defparam \mem[0][102] .is_wysiwyg = "true";
defparam \mem[0][102] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!in_ready_hold),
	.datab(!mem_used_1),
	.datac(!in_data_reg_60),
	.datad(!out_valid_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h0004000400040004;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h0202020202020202;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'h5545331355453313;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][117] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][117]~q ),
	.prn(vcc));
defparam \mem[1][117] .is_wysiwyg = "true";
defparam \mem[1][117] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!nxt_out_eop),
	.datac(!\mem[1][117]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!last_packet_beat),
	.datac(!read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hAEAEAEAEAEAEAEAE;
defparam \always0~0 .shared_arith = "off";

dffeas \mem[1][60] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][60]~q ),
	.prn(vcc));
defparam \mem[1][60] .is_wysiwyg = "true";
defparam \mem[1][60] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!mem_used_1),
	.datab(!in_data_reg_60),
	.datac(!\mem[1][60]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h2727272727272727;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!mem_used_0),
	.datac(!last_packet_beat),
	.datad(!read),
	.datae(!write1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h3313FFFF3313FFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem[1][69] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][69]~q ),
	.prn(vcc));
defparam \mem[1][69] .is_wysiwyg = "true";
defparam \mem[1][69] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!\mem[1][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h0257025702570257;
defparam \mem~2 .shared_arith = "off";

dffeas \mem[1][68] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][68]~q ),
	.prn(vcc));
defparam \mem[1][68] .is_wysiwyg = "true";
defparam \mem[1][68] .power_up = "low";

cyclonev_lcell_comb \mem~3 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\mem[1][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~3 .extended_lut = "off";
defparam \mem~3 .lut_mask = 64'h0257025702570257;
defparam \mem~3 .shared_arith = "off";

dffeas \mem[1][67] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][67]~q ),
	.prn(vcc));
defparam \mem[1][67] .is_wysiwyg = "true";
defparam \mem[1][67] .power_up = "low";

cyclonev_lcell_comb \mem~4 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!\mem[1][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~4 .extended_lut = "off";
defparam \mem~4 .lut_mask = 64'h0257025702570257;
defparam \mem~4 .shared_arith = "off";

dffeas \mem[1][66] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][66]~q ),
	.prn(vcc));
defparam \mem[1][66] .is_wysiwyg = "true";
defparam \mem[1][66] .power_up = "low";

cyclonev_lcell_comb \mem~5 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\mem[1][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~5 .extended_lut = "off";
defparam \mem~5 .lut_mask = 64'h0257025702570257;
defparam \mem~5 .shared_arith = "off";

dffeas \mem[1][65] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][65]~q ),
	.prn(vcc));
defparam \mem[1][65] .is_wysiwyg = "true";
defparam \mem[1][65] .power_up = "low";

cyclonev_lcell_comb \mem~6 (
	.dataa(!mem_used_1),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(!out_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(!\mem[1][65]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~6 .extended_lut = "off";
defparam \mem~6 .lut_mask = 64'h082A5D7F082A5D7F;
defparam \mem~6 .shared_arith = "off";

dffeas \mem[1][92] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][92]~q ),
	.prn(vcc));
defparam \mem[1][92] .is_wysiwyg = "true";
defparam \mem[1][92] .power_up = "low";

cyclonev_lcell_comb \mem~7 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][92]~q ),
	.datac(!in_data_reg_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~7 .extended_lut = "off";
defparam \mem~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~7 .shared_arith = "off";

dffeas \mem[1][93] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][93]~q ),
	.prn(vcc));
defparam \mem[1][93] .is_wysiwyg = "true";
defparam \mem[1][93] .power_up = "low";

cyclonev_lcell_comb \mem~8 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][93]~q ),
	.datac(!in_data_reg_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~8 .extended_lut = "off";
defparam \mem~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~8 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~9 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][94]~q ),
	.datac(!in_data_reg_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~9 .extended_lut = "off";
defparam \mem~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~9 .shared_arith = "off";

dffeas \mem[1][95] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][95]~q ),
	.prn(vcc));
defparam \mem[1][95] .is_wysiwyg = "true";
defparam \mem[1][95] .power_up = "low";

cyclonev_lcell_comb \mem~10 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][95]~q ),
	.datac(!in_data_reg_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~10 .extended_lut = "off";
defparam \mem~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~10 .shared_arith = "off";

dffeas \mem[1][96] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][96]~q ),
	.prn(vcc));
defparam \mem[1][96] .is_wysiwyg = "true";
defparam \mem[1][96] .power_up = "low";

cyclonev_lcell_comb \mem~11 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][96]~q ),
	.datac(!in_data_reg_96),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~11 .extended_lut = "off";
defparam \mem~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~11 .shared_arith = "off";

dffeas \mem[1][97] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][97]~q ),
	.prn(vcc));
defparam \mem[1][97] .is_wysiwyg = "true";
defparam \mem[1][97] .power_up = "low";

cyclonev_lcell_comb \mem~12 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][97]~q ),
	.datac(!in_data_reg_97),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~12 .extended_lut = "off";
defparam \mem~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~12 .shared_arith = "off";

dffeas \mem[1][98] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][98]~q ),
	.prn(vcc));
defparam \mem[1][98] .is_wysiwyg = "true";
defparam \mem[1][98] .power_up = "low";

cyclonev_lcell_comb \mem~13 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][98]~q ),
	.datac(!in_data_reg_98),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~13 .extended_lut = "off";
defparam \mem~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~13 .shared_arith = "off";

dffeas \mem[1][99] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][99]~q ),
	.prn(vcc));
defparam \mem[1][99] .is_wysiwyg = "true";
defparam \mem[1][99] .power_up = "low";

cyclonev_lcell_comb \mem~14 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][99]~q ),
	.datac(!in_data_reg_99),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~14 .extended_lut = "off";
defparam \mem~14 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~14 .shared_arith = "off";

dffeas \mem[1][100] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][100]~q ),
	.prn(vcc));
defparam \mem[1][100] .is_wysiwyg = "true";
defparam \mem[1][100] .power_up = "low";

cyclonev_lcell_comb \mem~15 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][100]~q ),
	.datac(!in_data_reg_100),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~15 .extended_lut = "off";
defparam \mem~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~15 .shared_arith = "off";

dffeas \mem[1][101] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][101]~q ),
	.prn(vcc));
defparam \mem[1][101] .is_wysiwyg = "true";
defparam \mem[1][101] .power_up = "low";

cyclonev_lcell_comb \mem~16 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][101]~q ),
	.datac(!in_data_reg_101),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~16 .extended_lut = "off";
defparam \mem~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~16 .shared_arith = "off";

dffeas \mem[1][102] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][102]~q ),
	.prn(vcc));
defparam \mem[1][102] .is_wysiwyg = "true";
defparam \mem[1][102] .power_up = "low";

cyclonev_lcell_comb \mem~17 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][102]~q ),
	.datac(!in_data_reg_102),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~17 .extended_lut = "off";
defparam \mem~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~17 .shared_arith = "off";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

cyclonev_lcell_comb \mem~18 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][103]~q ),
	.datac(!in_data_reg_103),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~18 .extended_lut = "off";
defparam \mem~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem~18 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_axi_master_ni (
	h2f_lw_AWVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_WVALID_0,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWADDR_15,
	h2f_lw_AWADDR_16,
	h2f_lw_AWADDR_17,
	h2f_lw_AWADDR_18,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_0,
	h2f_lw_AWLEN_1,
	h2f_lw_AWLEN_2,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	address_burst_7,
	address_burst_6,
	address_burst_9,
	address_burst_8,
	address_burst_11,
	address_burst_10,
	address_burst_15,
	address_burst_14,
	address_burst_13,
	address_burst_12,
	Add5,
	Add51,
	write_addr_data_both_valid1,
	sop_enable1,
	address_burst_5,
	address_burst_4,
	out_data_18,
	out_data_17,
	out_data_16,
	nonposted_cmd_accepted,
	Decoder1,
	Add2,
	Add21,
	Add22,
	altera_reset_synchronizer_int_chain_out,
	burst_bytecount_6,
	write_cp_data_69,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_2,
	write_cp_data_65,
	Selector3,
	Selector10,
	Selector101,
	base_address_3,
	Selector4,
	Selector11,
	base_address_2,
	Selector5,
	Add3,
	Selector12,
	out_data_1,
	Decoder11,
	out_data_0,
	Selector6,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_WVALID_0;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWADDR_15;
input 	h2f_lw_AWADDR_16;
input 	h2f_lw_AWADDR_17;
input 	h2f_lw_AWADDR_18;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_0;
input 	h2f_lw_AWLEN_1;
input 	h2f_lw_AWLEN_2;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
output 	address_burst_7;
output 	address_burst_6;
output 	address_burst_9;
output 	address_burst_8;
output 	address_burst_11;
output 	address_burst_10;
output 	address_burst_15;
output 	address_burst_14;
output 	address_burst_13;
output 	address_burst_12;
output 	Add5;
output 	Add51;
output 	write_addr_data_both_valid1;
output 	sop_enable1;
output 	address_burst_5;
output 	address_burst_4;
output 	out_data_18;
output 	out_data_17;
output 	out_data_16;
input 	nonposted_cmd_accepted;
output 	Decoder1;
output 	Add2;
output 	Add21;
output 	Add22;
input 	altera_reset_synchronizer_int_chain_out;
output 	burst_bytecount_6;
output 	write_cp_data_69;
output 	burst_bytecount_5;
output 	write_cp_data_68;
output 	burst_bytecount_4;
output 	write_cp_data_67;
output 	burst_bytecount_3;
output 	write_cp_data_66;
output 	burst_bytecount_2;
output 	write_cp_data_65;
output 	Selector3;
output 	Selector10;
output 	Selector101;
output 	base_address_3;
output 	Selector4;
output 	Selector11;
output 	base_address_2;
output 	Selector5;
output 	Add3;
output 	Selector12;
output 	out_data_1;
output 	Decoder11;
output 	out_data_0;
output 	Selector6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \LessThan14~0_combout ;
wire \align_address_to_size|Selector17~0_combout ;
wire \align_address_to_size|Decoder0~4_combout ;
wire \align_address_to_size|Decoder0~5_combout ;
wire \align_address_to_size|Decoder0~6_combout ;
wire \align_address_to_size|Decoder0~7_combout ;
wire \Add5~10 ;
wire \Add5~14 ;
wire \Decoder1~3_combout ;
wire \sop_enable~0_combout ;
wire \Add7~0_combout ;
wire \Add0~0_combout ;
wire \Add7~1_combout ;
wire \Add7~2_combout ;
wire \Add7~3_combout ;
wire \Add4~14 ;
wire \Add4~10 ;
wire \Add4~6 ;
wire \Add4~1_sumout ;
wire \Add3~0_combout ;
wire \Decoder1~1_combout ;
wire \Decoder1~2_combout ;
wire \Add5~6 ;
wire \Add5~1_sumout ;
wire \log2ceil~0_combout ;
wire \Add1~0_combout ;
wire \Add1~1_combout ;
wire \Selector4~0_combout ;
wire \Add4~5_sumout ;
wire \Add3~1_combout ;
wire \Add3~2_combout ;
wire \Add5~5_sumout ;
wire \Selector11~0_combout ;
wire \Add4~9_sumout ;
wire \Selector5~0_combout ;
wire \Add4~13_sumout ;


terminal_qsys_altera_merlin_address_alignment align_address_to_size(
	.h2f_lw_AWADDR_0(h2f_lw_AWADDR_0),
	.h2f_lw_AWADDR_1(h2f_lw_AWADDR_1),
	.h2f_lw_AWADDR_2(h2f_lw_AWADDR_2),
	.h2f_lw_AWADDR_3(h2f_lw_AWADDR_3),
	.h2f_lw_AWADDR_4(h2f_lw_AWADDR_4),
	.h2f_lw_AWADDR_5(h2f_lw_AWADDR_5),
	.h2f_lw_AWADDR_6(h2f_lw_AWADDR_6),
	.h2f_lw_AWADDR_7(h2f_lw_AWADDR_7),
	.h2f_lw_AWADDR_8(h2f_lw_AWADDR_8),
	.h2f_lw_AWADDR_9(h2f_lw_AWADDR_9),
	.h2f_lw_AWADDR_10(h2f_lw_AWADDR_10),
	.h2f_lw_AWADDR_11(h2f_lw_AWADDR_11),
	.h2f_lw_AWADDR_12(h2f_lw_AWADDR_12),
	.h2f_lw_AWADDR_13(h2f_lw_AWADDR_13),
	.h2f_lw_AWADDR_14(h2f_lw_AWADDR_14),
	.h2f_lw_AWADDR_15(h2f_lw_AWADDR_15),
	.h2f_lw_AWADDR_16(h2f_lw_AWADDR_16),
	.h2f_lw_AWADDR_17(h2f_lw_AWADDR_17),
	.h2f_lw_AWADDR_18(h2f_lw_AWADDR_18),
	.h2f_lw_AWBURST_0(h2f_lw_AWBURST_0),
	.h2f_lw_AWBURST_1(h2f_lw_AWBURST_1),
	.h2f_lw_AWLEN_3(h2f_lw_AWLEN_3),
	.h2f_lw_AWSIZE_0(h2f_lw_AWSIZE_0),
	.h2f_lw_AWSIZE_1(h2f_lw_AWSIZE_1),
	.h2f_lw_AWSIZE_2(h2f_lw_AWSIZE_2),
	.address_burst_7(address_burst_7),
	.address_burst_6(address_burst_6),
	.address_burst_9(address_burst_9),
	.address_burst_8(address_burst_8),
	.address_burst_11(address_burst_11),
	.address_burst_10(address_burst_10),
	.address_burst_15(address_burst_15),
	.address_burst_14(address_burst_14),
	.address_burst_13(address_burst_13),
	.address_burst_12(address_burst_12),
	.sop_enable(sop_enable1),
	.address_burst_5(address_burst_5),
	.address_burst_4(address_burst_4),
	.out_data_18(out_data_18),
	.out_data_17(out_data_17),
	.out_data_16(out_data_16),
	.nonposted_cmd_accepted(nonposted_cmd_accepted),
	.reset(altera_reset_synchronizer_int_chain_out),
	.log2ceil(\log2ceil~0_combout ),
	.Add1(\Add1~0_combout ),
	.Add11(\Add1~1_combout ),
	.LessThan14(\LessThan14~0_combout ),
	.Selector17(\align_address_to_size|Selector17~0_combout ),
	.base_address_3(base_address_3),
	.Selector4(\Selector4~0_combout ),
	.base_address_2(base_address_2),
	.Decoder0(\align_address_to_size|Decoder0~4_combout ),
	.Decoder01(\align_address_to_size|Decoder0~5_combout ),
	.Decoder02(\align_address_to_size|Decoder0~6_combout ),
	.Selector5(\Selector5~0_combout ),
	.out_data_1(out_data_1),
	.Decoder03(\align_address_to_size|Decoder0~7_combout ),
	.out_data_0(out_data_0),
	.clk(clk_clk));

cyclonev_lcell_comb \LessThan14~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan14~0 .extended_lut = "off";
defparam \LessThan14~0 .lut_mask = 64'hE8A0A080A0808000;
defparam \LessThan14~0 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add5),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h00000000000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Decoder11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add51),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h00000000000000FF;
defparam \Add5~13 .shared_arith = "off";

cyclonev_lcell_comb write_addr_data_both_valid(
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_addr_data_both_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam write_addr_data_both_valid.extended_lut = "off";
defparam write_addr_data_both_valid.lut_mask = 64'h1111111111111111;
defparam write_addr_data_both_valid.shared_arith = "off";

dffeas sop_enable(
	.clk(clk_clk),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(sop_enable1),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

cyclonev_lcell_comb \Decoder1~0 (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~0 .extended_lut = "off";
defparam \Decoder1~0 .lut_mask = 64'h8888888888888888;
defparam \Decoder1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \Add2~0 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h01FE01FE01FE01FE;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~2 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~2 .extended_lut = "off";
defparam \Add2~2 .lut_mask = 64'h0001000100010001;
defparam \Add2~2 .shared_arith = "off";

dffeas \burst_bytecount[6] (
	.clk(clk_clk),
	.d(\Add7~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_6),
	.prn(vcc));
defparam \burst_bytecount[6] .is_wysiwyg = "true";
defparam \burst_bytecount[6] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[69]~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_6),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_69),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[69]~0 .extended_lut = "off";
defparam \write_cp_data[69]~0 .lut_mask = 64'h0347034703470347;
defparam \write_cp_data[69]~0 .shared_arith = "off";

dffeas \burst_bytecount[5] (
	.clk(clk_clk),
	.d(\Add7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_5),
	.prn(vcc));
defparam \burst_bytecount[5] .is_wysiwyg = "true";
defparam \burst_bytecount[5] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[68]~1 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!sop_enable1),
	.datac(!\Add0~0_combout ),
	.datad(!burst_bytecount_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_68),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[68]~1 .extended_lut = "off";
defparam \write_cp_data[68]~1 .lut_mask = 64'h487B487B487B487B;
defparam \write_cp_data[68]~1 .shared_arith = "off";

dffeas \burst_bytecount[4] (
	.clk(clk_clk),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_4),
	.prn(vcc));
defparam \burst_bytecount[4] .is_wysiwyg = "true";
defparam \burst_bytecount[4] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[67]~2 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!sop_enable1),
	.datae(!burst_bytecount_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_67),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[67]~2 .extended_lut = "off";
defparam \write_cp_data[67]~2 .lut_mask = 64'h1E001EFF1E001EFF;
defparam \write_cp_data[67]~2 .shared_arith = "off";

dffeas \burst_bytecount[3] (
	.clk(clk_clk),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_3),
	.prn(vcc));
defparam \burst_bytecount[3] .is_wysiwyg = "true";
defparam \burst_bytecount[3] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[66]~3 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!sop_enable1),
	.datad(!burst_bytecount_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_66),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[66]~3 .extended_lut = "off";
defparam \write_cp_data[66]~3 .lut_mask = 64'h606F606F606F606F;
defparam \write_cp_data[66]~3 .shared_arith = "off";

dffeas \burst_bytecount[2] (
	.clk(clk_clk),
	.d(write_cp_data_65),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(burst_bytecount_2),
	.prn(vcc));
defparam \burst_bytecount[2] .is_wysiwyg = "true";
defparam \burst_bytecount[2] .power_up = "low";

cyclonev_lcell_comb \write_cp_data[65]~4 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!sop_enable1),
	.datac(!burst_bytecount_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_cp_data_65),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_cp_data[65]~4 .extended_lut = "off";
defparam \write_cp_data[65]~4 .lut_mask = 64'h7474747474747474;
defparam \write_cp_data[65]~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add4~1_sumout ),
	.datad(!\align_address_to_size|Selector17~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h80A280A280A280A2;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\Add3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h8080808080808080;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Add5~1_sumout ),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector101),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h7F5D7F5D7F5D7F5D;
defparam \Selector10~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Selector4~0_combout ),
	.datad(!\Add4~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'h8A028A028A028A02;
defparam \Selector4~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~1 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Add3~1_combout ),
	.datad(!\Add3~2_combout ),
	.datae(!\Add5~5_sumout ),
	.dataf(!\Selector11~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~1 .extended_lut = "off";
defparam \Selector11~1 .lut_mask = 64'h5777DFFF7777FFFF;
defparam \Selector11~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add4~9_sumout ),
	.datad(!\Selector5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'h80A280A280A280A2;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~3 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Add3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~3 .extended_lut = "off";
defparam \Add3~3 .lut_mask = 64'h3F007000C0FF8FFF;
defparam \Add3~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector12~0 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!\Add3~1_combout ),
	.datad(!\Add3~2_combout ),
	.datae(!Add3),
	.dataf(!Add5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "off";
defparam \Selector12~0 .lut_mask = 64'h57777777DFFFFFFF;
defparam \Selector12~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~4 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~4 .extended_lut = "off";
defparam \Decoder1~4 .lut_mask = 64'h8080808080808080;
defparam \Decoder1~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add1~1_combout ),
	.datad(!\Add4~13_sumout ),
	.datae(!\Selector5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h8800A8208800A820;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~3 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~3 .extended_lut = "off";
defparam \Decoder1~3 .lut_mask = 64'h4040404040404040;
defparam \Decoder1~3 .shared_arith = "off";

cyclonev_lcell_comb \sop_enable~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_enable~0 .extended_lut = "off";
defparam \sop_enable~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sop_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!write_cp_data_69),
	.datab(!write_cp_data_68),
	.datac(!write_cp_data_66),
	.datad(!write_cp_data_65),
	.datae(!write_cp_data_67),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h5595555555955555;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h0101010101010101;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!write_cp_data_68),
	.datab(!write_cp_data_66),
	.datac(!write_cp_data_65),
	.datad(!write_cp_data_67),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h5955595559555955;
defparam \Add7~1 .shared_arith = "off";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!write_cp_data_66),
	.datab(!write_cp_data_65),
	.datac(!write_cp_data_67),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h2D2D2D2D2D2D2D2D;
defparam \Add7~2 .shared_arith = "off";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!write_cp_data_66),
	.datab(!write_cp_data_65),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h6666666666666666;
defparam \Add7~3 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\align_address_to_size|Decoder0~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~0 .extended_lut = "off";
defparam \Add3~0 .lut_mask = 64'h00000F003F007F00;
defparam \Add3~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~1 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~1 .extended_lut = "off";
defparam \Decoder1~1 .lut_mask = 64'h1010101010101010;
defparam \Decoder1~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder1~2 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_ARSIZE_1),
	.datac(!h2f_lw_ARSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder1~2 .extended_lut = "off";
defparam \Decoder1~2 .lut_mask = 64'h2020202020202020;
defparam \Decoder1~2 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~5_sumout ),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h00000000000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Decoder1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~1_sumout ),
	.cout(),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h00000000000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \log2ceil~0 (
	.dataa(!h2f_lw_AWLEN_1),
	.datab(!h2f_lw_AWLEN_2),
	.datac(!h2f_lw_AWLEN_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\log2ceil~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \log2ceil~0 .extended_lut = "off";
defparam \log2ceil~0 .lut_mask = 64'h7070707070707070;
defparam \log2ceil~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h00004F0000004F00;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!h2f_lw_AWLEN_0),
	.datab(!h2f_lw_AWLEN_1),
	.datac(!h2f_lw_AWLEN_2),
	.datad(!h2f_lw_AWLEN_3),
	.datae(!h2f_lw_AWSIZE_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4F00B0FF4F00B0FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'hA080800080000000;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\Add3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h1717171717171717;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add3~2 (
	.dataa(!h2f_lw_ARLEN_3),
	.datab(!h2f_lw_ARSIZE_2),
	.datac(!\Add3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add3~2 .extended_lut = "off";
defparam \Add3~2 .lut_mask = 64'h6969696969696969;
defparam \Add3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(!h2f_lw_ARSIZE_0),
	.dataf(!h2f_lw_ARSIZE_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h0F003000400080FF;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!\log2ceil~0_combout ),
	.datae(!\Add1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h8000000080000000;
defparam \Selector5~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_address_alignment (
	h2f_lw_AWADDR_0,
	h2f_lw_AWADDR_1,
	h2f_lw_AWADDR_2,
	h2f_lw_AWADDR_3,
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWADDR_15,
	h2f_lw_AWADDR_16,
	h2f_lw_AWADDR_17,
	h2f_lw_AWADDR_18,
	h2f_lw_AWBURST_0,
	h2f_lw_AWBURST_1,
	h2f_lw_AWLEN_3,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	address_burst_7,
	address_burst_6,
	address_burst_9,
	address_burst_8,
	address_burst_11,
	address_burst_10,
	address_burst_15,
	address_burst_14,
	address_burst_13,
	address_burst_12,
	sop_enable,
	address_burst_5,
	address_burst_4,
	out_data_18,
	out_data_17,
	out_data_16,
	nonposted_cmd_accepted,
	reset,
	log2ceil,
	Add1,
	Add11,
	LessThan14,
	Selector17,
	base_address_3,
	Selector4,
	base_address_2,
	Decoder0,
	Decoder01,
	Decoder02,
	Selector5,
	out_data_1,
	Decoder03,
	out_data_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_0;
input 	h2f_lw_AWADDR_1;
input 	h2f_lw_AWADDR_2;
input 	h2f_lw_AWADDR_3;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWADDR_15;
input 	h2f_lw_AWADDR_16;
input 	h2f_lw_AWADDR_17;
input 	h2f_lw_AWADDR_18;
input 	h2f_lw_AWBURST_0;
input 	h2f_lw_AWBURST_1;
input 	h2f_lw_AWLEN_3;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
output 	address_burst_7;
output 	address_burst_6;
output 	address_burst_9;
output 	address_burst_8;
output 	address_burst_11;
output 	address_burst_10;
output 	address_burst_15;
output 	address_burst_14;
output 	address_burst_13;
output 	address_burst_12;
input 	sop_enable;
output 	address_burst_5;
output 	address_burst_4;
output 	out_data_18;
output 	out_data_17;
output 	out_data_16;
input 	nonposted_cmd_accepted;
input 	reset;
input 	log2ceil;
input 	Add1;
input 	Add11;
input 	LessThan14;
output 	Selector17;
output 	base_address_3;
input 	Selector4;
output 	base_address_2;
output 	Decoder0;
output 	Decoder01;
output 	Decoder02;
input 	Selector5;
output 	out_data_1;
output 	Decoder03;
output 	out_data_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Decoder0~2_combout ;
wire \Decoder0~3_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \Add0~73_sumout ;
wire \Add1~21_sumout ;
wire \Selector20~0_combout ;
wire \address_burst[0]~q ;
wire \Add1~22 ;
wire \Add1~17_sumout ;
wire \aligned_address_bits[1]~combout ;
wire \Add0~74 ;
wire \Add0~69_sumout ;
wire \Selector19~0_combout ;
wire \address_burst[1]~q ;
wire \Add1~18 ;
wire \Add1~13_sumout ;
wire \Add0~70 ;
wire \Add0~65_sumout ;
wire \Selector18~0_combout ;
wire \address_burst[2]~q ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \Add0~66 ;
wire \Add0~61_sumout ;
wire \Selector17~1_combout ;
wire \address_burst[3]~q ;
wire \Add0~62 ;
wire \Add0~6 ;
wire \Add0~2 ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \out_data[7]~5_combout ;
wire \Add0~13_sumout ;
wire \out_data[6]~6_combout ;
wire \Add0~10 ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \out_data[9]~7_combout ;
wire \Add0~21_sumout ;
wire \out_data[8]~8_combout ;
wire \Add0~18 ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \out_data[11]~9_combout ;
wire \Add0~29_sumout ;
wire \out_data[10]~10_combout ;
wire \Add0~26 ;
wire \Add0~46 ;
wire \Add0~42 ;
wire \Add0~38 ;
wire \Add0~33_sumout ;
wire \out_data[15]~11_combout ;
wire \Add0~37_sumout ;
wire \out_data[14]~12_combout ;
wire \Add0~41_sumout ;
wire \out_data[13]~13_combout ;
wire \Add0~45_sumout ;
wire \out_data[12]~14_combout ;
wire \out_data[5]~3_combout ;
wire \Add1~10 ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \Selector15~0_combout ;
wire \Add0~1_sumout ;
wire \Selector15~1_combout ;
wire \out_data[4]~4_combout ;
wire \Add1~5_sumout ;
wire \Add0~5_sumout ;
wire \Selector16~0_combout ;
wire \Add0~34 ;
wire \Add0~57_sumout ;
wire \address_burst[16]~q ;
wire \Add0~58 ;
wire \Add0~53_sumout ;
wire \address_burst[17]~q ;
wire \Add0~54 ;
wire \Add0~49_sumout ;
wire \address_burst[18]~q ;


dffeas \address_burst[7] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(\out_data[7]~5_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_7),
	.prn(vcc));
defparam \address_burst[7] .is_wysiwyg = "true";
defparam \address_burst[7] .power_up = "low";

dffeas \address_burst[6] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(\out_data[6]~6_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_6),
	.prn(vcc));
defparam \address_burst[6] .is_wysiwyg = "true";
defparam \address_burst[6] .power_up = "low";

dffeas \address_burst[9] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(\out_data[9]~7_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_9),
	.prn(vcc));
defparam \address_burst[9] .is_wysiwyg = "true";
defparam \address_burst[9] .power_up = "low";

dffeas \address_burst[8] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(\out_data[8]~8_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_8),
	.prn(vcc));
defparam \address_burst[8] .is_wysiwyg = "true";
defparam \address_burst[8] .power_up = "low";

dffeas \address_burst[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(\out_data[11]~9_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_11),
	.prn(vcc));
defparam \address_burst[11] .is_wysiwyg = "true";
defparam \address_burst[11] .power_up = "low";

dffeas \address_burst[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(\out_data[10]~10_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_10),
	.prn(vcc));
defparam \address_burst[10] .is_wysiwyg = "true";
defparam \address_burst[10] .power_up = "low";

dffeas \address_burst[15] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(\out_data[15]~11_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_15),
	.prn(vcc));
defparam \address_burst[15] .is_wysiwyg = "true";
defparam \address_burst[15] .power_up = "low";

dffeas \address_burst[14] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(\out_data[14]~12_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_14),
	.prn(vcc));
defparam \address_burst[14] .is_wysiwyg = "true";
defparam \address_burst[14] .power_up = "low";

dffeas \address_burst[13] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(\out_data[13]~13_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_13),
	.prn(vcc));
defparam \address_burst[13] .is_wysiwyg = "true";
defparam \address_burst[13] .power_up = "low";

dffeas \address_burst[12] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(\out_data[12]~14_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_12),
	.prn(vcc));
defparam \address_burst[12] .is_wysiwyg = "true";
defparam \address_burst[12] .power_up = "low";

dffeas \address_burst[5] (
	.clk(clk),
	.d(\Selector15~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_5),
	.prn(vcc));
defparam \address_burst[5] .is_wysiwyg = "true";
defparam \address_burst[5] .power_up = "low";

dffeas \address_burst[4] (
	.clk(clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(address_burst_4),
	.prn(vcc));
defparam \address_burst[4] .is_wysiwyg = "true";
defparam \address_burst[4] .power_up = "low";

cyclonev_lcell_comb \out_data[18]~0 (
	.dataa(!h2f_lw_AWADDR_18),
	.datab(!sop_enable),
	.datac(!\address_burst[18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[18]~0 .extended_lut = "off";
defparam \out_data[18]~0 .lut_mask = 64'h4747474747474747;
defparam \out_data[18]~0 .shared_arith = "off";

cyclonev_lcell_comb \out_data[17]~1 (
	.dataa(!h2f_lw_AWADDR_17),
	.datab(!sop_enable),
	.datac(!\address_burst[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[17]~1 .extended_lut = "off";
defparam \out_data[17]~1 .lut_mask = 64'h4747474747474747;
defparam \out_data[17]~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[16]~2 (
	.dataa(!h2f_lw_AWADDR_16),
	.datab(!sop_enable),
	.datac(!\address_burst[16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[16]~2 .extended_lut = "off";
defparam \out_data[16]~2 .lut_mask = 64'h4747474747474747;
defparam \out_data[16]~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!log2ceil),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector17),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'hA0808000A0808000;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \base_address[3]~0 (
	.dataa(!h2f_lw_AWADDR_3),
	.datab(!sop_enable),
	.datac(!\address_burst[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[3]~0 .extended_lut = "off";
defparam \base_address[3]~0 .lut_mask = 64'h4747474747474747;
defparam \base_address[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \base_address[2]~1 (
	.dataa(!h2f_lw_AWADDR_2),
	.datab(!sop_enable),
	.datac(!\address_burst[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(base_address_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \base_address[2]~1 .extended_lut = "off";
defparam \base_address[2]~1 .lut_mask = 64'h4747474747474747;
defparam \base_address[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~4 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~4 .extended_lut = "off";
defparam \Decoder0~4 .lut_mask = 64'h1010101010101010;
defparam \Decoder0~4 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~5 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~5 .extended_lut = "off";
defparam \Decoder0~5 .lut_mask = 64'h2020202020202020;
defparam \Decoder0~5 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~6 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder02),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~6 .extended_lut = "off";
defparam \Decoder0~6 .lut_mask = 64'h4040404040404040;
defparam \Decoder0~6 .shared_arith = "off";

cyclonev_lcell_comb \out_data[1]~15 (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!sop_enable),
	.datac(!\address_burst[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[1]~15 .extended_lut = "off";
defparam \out_data[1]~15 .lut_mask = 64'h4747474747474747;
defparam \out_data[1]~15 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~7 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Decoder03),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~7 .extended_lut = "off";
defparam \Decoder0~7 .lut_mask = 64'h8080808080808080;
defparam \Decoder0~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[0]~16 (
	.dataa(!h2f_lw_AWADDR_0),
	.datab(!sop_enable),
	.datac(!\address_burst[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(out_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[0]~16 .extended_lut = "off";
defparam \out_data[0]~16 .lut_mask = 64'h4747474747474747;
defparam \out_data[0]~16 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'h0101010101010101;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~3 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~3 .extended_lut = "off";
defparam \Decoder0~3 .lut_mask = 64'h0202020202020202;
defparam \Decoder0~3 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h0404040404040404;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!h2f_lw_AWSIZE_0),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'h0808080808080808;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~73 (
	.dataa(!sop_enable),
	.datab(!\address_burst[0]~q ),
	.datac(!h2f_lw_AWADDR_0),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!Decoder03),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h0000EEE4000000FF;
defparam \Add0~73 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[0]~q ),
	.datad(!Decoder03),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Selector20~0 (
	.dataa(!Add11),
	.datab(!out_data_0),
	.datac(!\Add0~73_sumout ),
	.datad(!\Add1~21_sumout ),
	.datae(!h2f_lw_AWBURST_0),
	.dataf(!h2f_lw_AWBURST_1),
	.datag(!Selector5),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "on";
defparam \Selector20~0 .lut_mask = 64'h33330F0F02F70F0F;
defparam \Selector20~0 .shared_arith = "off";

dffeas \address_burst[0] (
	.clk(clk),
	.d(\Selector20~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[0]~q ),
	.prn(vcc));
defparam \address_burst[0] .is_wysiwyg = "true";
defparam \address_burst[0] .power_up = "low";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!h2f_lw_AWADDR_1),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FA50000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \aligned_address_bits[1] (
	.dataa(!h2f_lw_AWADDR_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aligned_address_bits[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aligned_address_bits[1] .extended_lut = "off";
defparam \aligned_address_bits[1] .lut_mask = 64'h4040404040404040;
defparam \aligned_address_bits[1] .shared_arith = "off";

cyclonev_lcell_comb \Add0~69 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!\address_burst[1]~q ),
	.datad(!Decoder02),
	.datae(gnd),
	.dataf(!\aligned_address_bits[1]~combout ),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h0000FA50000000FF;
defparam \Add0~69 .shared_arith = "off";

cyclonev_lcell_comb \Selector19~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\Add1~17_sumout ),
	.datad(!\Add0~69_sumout ),
	.datae(!Selector5),
	.dataf(!out_data_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h025700558ADFAAFF;
defparam \Selector19~0 .shared_arith = "off";

dffeas \address_burst[1] (
	.clk(clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[1]~q ),
	.prn(vcc));
defparam \address_burst[1] .is_wysiwyg = "true";
defparam \address_burst[1] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_2),
	.datad(!Decoder01),
	.datae(gnd),
	.dataf(!\address_burst[2]~q ),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~65 .shared_arith = "off";

cyclonev_lcell_comb \Selector18~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Selector4),
	.datad(!base_address_2),
	.datae(!\Add1~13_sumout ),
	.dataf(!\Add0~65_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector18~0 .extended_lut = "off";
defparam \Selector18~0 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector18~0 .shared_arith = "off";

dffeas \address_burst[2] (
	.clk(clk),
	.d(\Selector18~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[2]~q ),
	.prn(vcc));
defparam \address_burst[2] .is_wysiwyg = "true";
defparam \address_burst[2] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_3),
	.datad(!Decoder0),
	.datae(gnd),
	.dataf(!\address_burst[3]~q ),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Selector17~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!Selector17),
	.datad(!base_address_3),
	.datae(!\Add1~9_sumout ),
	.dataf(!\Add0~61_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~1 .extended_lut = "off";
defparam \Selector17~1 .lut_mask = 64'h008A20AA55DF75FF;
defparam \Selector17~1 .shared_arith = "off";

dffeas \address_burst[3] (
	.clk(clk),
	.d(\Selector17~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[3]~q ),
	.prn(vcc));
defparam \address_burst[3] .is_wysiwyg = "true";
defparam \address_burst[3] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!address_burst_4),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_5),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!address_burst_5),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_6),
	.datad(!\Decoder0~3_combout ),
	.datae(gnd),
	.dataf(!address_burst_6),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_7),
	.datad(!\Decoder0~2_combout ),
	.datae(gnd),
	.dataf(!address_burst_7),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \out_data[7]~5 (
	.dataa(!h2f_lw_AWADDR_7),
	.datab(!sop_enable),
	.datac(!address_burst_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[7]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[7]~5 .extended_lut = "off";
defparam \out_data[7]~5 .lut_mask = 64'h4747474747474747;
defparam \out_data[7]~5 .shared_arith = "off";

cyclonev_lcell_comb \out_data[6]~6 (
	.dataa(!h2f_lw_AWADDR_6),
	.datab(!sop_enable),
	.datac(!address_burst_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[6]~6 .extended_lut = "off";
defparam \out_data[6]~6 .lut_mask = 64'h4747474747474747;
defparam \out_data[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_8),
	.datad(!address_burst_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_9),
	.datad(!address_burst_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \out_data[9]~7 (
	.dataa(!h2f_lw_AWADDR_9),
	.datab(!sop_enable),
	.datac(!address_burst_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[9]~7 .extended_lut = "off";
defparam \out_data[9]~7 .lut_mask = 64'h4747474747474747;
defparam \out_data[9]~7 .shared_arith = "off";

cyclonev_lcell_comb \out_data[8]~8 (
	.dataa(!h2f_lw_AWADDR_8),
	.datab(!sop_enable),
	.datac(!address_burst_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[8]~8 .extended_lut = "off";
defparam \out_data[8]~8 .lut_mask = 64'h4747474747474747;
defparam \out_data[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_10),
	.datad(!address_burst_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_11),
	.datad(!address_burst_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \out_data[11]~9 (
	.dataa(!h2f_lw_AWADDR_11),
	.datab(!sop_enable),
	.datac(!address_burst_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[11]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[11]~9 .extended_lut = "off";
defparam \out_data[11]~9 .lut_mask = 64'h4747474747474747;
defparam \out_data[11]~9 .shared_arith = "off";

cyclonev_lcell_comb \out_data[10]~10 (
	.dataa(!h2f_lw_AWADDR_10),
	.datab(!sop_enable),
	.datac(!address_burst_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[10]~10 .extended_lut = "off";
defparam \out_data[10]~10 .lut_mask = 64'h4747474747474747;
defparam \out_data[10]~10 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_12),
	.datad(!address_burst_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_13),
	.datad(!address_burst_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_14),
	.datad(!address_burst_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_15),
	.datad(!address_burst_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \out_data[15]~11 (
	.dataa(!h2f_lw_AWADDR_15),
	.datab(!sop_enable),
	.datac(!address_burst_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[15]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[15]~11 .extended_lut = "off";
defparam \out_data[15]~11 .lut_mask = 64'h4747474747474747;
defparam \out_data[15]~11 .shared_arith = "off";

cyclonev_lcell_comb \out_data[14]~12 (
	.dataa(!h2f_lw_AWADDR_14),
	.datab(!sop_enable),
	.datac(!address_burst_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[14]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[14]~12 .extended_lut = "off";
defparam \out_data[14]~12 .lut_mask = 64'h4747474747474747;
defparam \out_data[14]~12 .shared_arith = "off";

cyclonev_lcell_comb \out_data[13]~13 (
	.dataa(!h2f_lw_AWADDR_13),
	.datab(!sop_enable),
	.datac(!address_burst_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[13]~13 .extended_lut = "off";
defparam \out_data[13]~13 .lut_mask = 64'h4747474747474747;
defparam \out_data[13]~13 .shared_arith = "off";

cyclonev_lcell_comb \out_data[12]~14 (
	.dataa(!h2f_lw_AWADDR_12),
	.datab(!sop_enable),
	.datac(!address_burst_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[12]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[12]~14 .extended_lut = "off";
defparam \out_data[12]~14 .lut_mask = 64'h4747474747474747;
defparam \out_data[12]~14 .shared_arith = "off";

cyclonev_lcell_comb \out_data[5]~3 (
	.dataa(!h2f_lw_AWADDR_5),
	.datab(!sop_enable),
	.datac(!address_burst_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[5]~3 .extended_lut = "off";
defparam \out_data[5]~3 .lut_mask = 64'h4747474747474747;
defparam \out_data[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_4),
	.datad(!\Decoder0~1_combout ),
	.datae(gnd),
	.dataf(!address_burst_4),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_5),
	.datad(!\Decoder0~0_combout ),
	.datae(gnd),
	.dataf(!address_burst_5),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000F5A0000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~0 (
	.dataa(!h2f_lw_AWLEN_3),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!h2f_lw_AWSIZE_2),
	.datad(!log2ceil),
	.datae(!Add1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'hE8A0A080E8A0A080;
defparam \Selector15~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector15~1 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\out_data[5]~3_combout ),
	.datad(!\Add1~1_sumout ),
	.datae(!\Selector15~0_combout ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~1 .extended_lut = "off";
defparam \Selector15~1 .lut_mask = 64'h082A0A0A5D7F5F5F;
defparam \Selector15~1 .shared_arith = "off";

cyclonev_lcell_comb \out_data[4]~4 (
	.dataa(!h2f_lw_AWADDR_4),
	.datab(!sop_enable),
	.datac(!address_burst_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_data[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_data[4]~4 .extended_lut = "off";
defparam \out_data[4]~4 .lut_mask = 64'h4747474747474747;
defparam \out_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector16~0 (
	.dataa(!h2f_lw_AWBURST_0),
	.datab(!h2f_lw_AWBURST_1),
	.datac(!\out_data[4]~4_combout ),
	.datad(!\Add1~5_sumout ),
	.datae(!LessThan14),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector16~0 .extended_lut = "off";
defparam \Selector16~0 .lut_mask = 64'h082A0A0A5D7F5F5F;
defparam \Selector16~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_16),
	.datad(!\address_burst[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~57 .shared_arith = "off";

dffeas \address_burst[16] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(out_data_16),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[16]~q ),
	.prn(vcc));
defparam \address_burst[16] .is_wysiwyg = "true";
defparam \address_burst[16] .power_up = "low";

cyclonev_lcell_comb \Add0~53 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_17),
	.datad(!\address_burst[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~53 .shared_arith = "off";

dffeas \address_burst[17] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(out_data_17),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[17]~q ),
	.prn(vcc));
defparam \address_burst[17] .is_wysiwyg = "true";
defparam \address_burst[17] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(!sop_enable),
	.datab(gnd),
	.datac(!h2f_lw_AWADDR_18),
	.datad(!\address_burst[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FFFF00000A5F;
defparam \Add0~49 .shared_arith = "off";

dffeas \address_burst[18] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(out_data_18),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(!h2f_lw_AWBURST_0),
	.ena(nonposted_cmd_accepted),
	.q(\address_burst[18]~q ),
	.prn(vcc));
defparam \address_burst[18] .is_wysiwyg = "true";
defparam \address_burst[18] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_burst_adapter (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	nxt_in_ready,
	saved_grant_1,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_ready_hold,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_59,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	Equal3,
	Equal4,
	saved_grant_0,
	in_data_reg_0,
	altera_reset_synchronizer_int_chain_out,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	Add2,
	Add21,
	Add22,
	src3_valid,
	src_valid,
	src_payload_0,
	nxt_out_eop,
	cp_ready,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	write_cp_data_69,
	write_cp_data_68,
	write_cp_data_67,
	write_cp_data_66,
	write_cp_data_65,
	WideNor0,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	src_payload,
	src_data_73,
	base_address_3,
	src_data_72,
	base_address_2,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	src_data_77,
	src_data_71,
	out_data_1,
	out_data_0,
	src_data_70,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
output 	nxt_in_ready;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_ready_hold;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_59;
input 	write;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	Equal3;
input 	Equal4;
input 	saved_grant_0;
output 	in_data_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	Add2;
input 	Add21;
input 	Add22;
input 	src3_valid;
input 	src_valid;
input 	src_payload_0;
output 	nxt_out_eop;
input 	cp_ready;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	write_cp_data_69;
input 	write_cp_data_68;
input 	write_cp_data_67;
input 	write_cp_data_66;
input 	write_cp_data_65;
input 	WideNor0;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	src_payload;
input 	src_data_73;
input 	base_address_3;
input 	src_data_72;
input 	base_address_2;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_100;
input 	src_data_101;
input 	src_data_102;
input 	src_data_103;
input 	src_data_77;
input 	src_data_71;
input 	out_data_1;
input 	out_data_0;
input 	src_data_70;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_adapter_13_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.nxt_in_ready(nxt_in_ready),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_103,src_data_102,src_data_101,src_data_100,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,src_data_77,gnd,gnd,gnd,
src_data_73,src_data_72,src_data_71,src_data_70,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,src_payload31,src_payload30,src_payload29,
src_payload28,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,src_payload10,
src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_ready_hold1(in_ready_hold),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_59(in_data_reg_59),
	.write(write),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal3(Equal3),
	.Equal4(Equal4),
	.in_data_reg_0(in_data_reg_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.src3_valid(src3_valid),
	.src_valid(src_valid),
	.sink0_endofpacket(src_payload_0),
	.nxt_out_eop(nxt_out_eop),
	.cp_ready(cp_ready),
	.in_data_reg_60(in_data_reg_60),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.write_cp_data_69(write_cp_data_69),
	.write_cp_data_68(write_cp_data_68),
	.write_cp_data_67(write_cp_data_67),
	.write_cp_data_66(write_cp_data_66),
	.write_cp_data_65(write_cp_data_65),
	.WideNor0(WideNor0),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_100(in_data_reg_100),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.base_address_3(base_address_3),
	.base_address_2(base_address_2),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_merlin_burst_adapter_13_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	nxt_in_ready,
	sink0_data,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_ready_hold1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_59,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	Equal3,
	Equal4,
	in_data_reg_0,
	altera_reset_synchronizer_int_chain_out,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	Add2,
	Add21,
	Add22,
	src3_valid,
	src_valid,
	sink0_endofpacket,
	nxt_out_eop,
	cp_ready,
	in_data_reg_60,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_6,
	write_cp_data_69,
	write_cp_data_68,
	write_cp_data_67,
	write_cp_data_66,
	write_cp_data_65,
	WideNor0,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	base_address_3,
	base_address_2,
	out_data_1,
	out_data_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
output 	nxt_in_ready;
input 	[115:0] sink0_data;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_ready_hold1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_59;
input 	write;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	Equal3;
input 	Equal4;
output 	in_data_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	Add2;
input 	Add21;
input 	Add22;
input 	src3_valid;
input 	src_valid;
input 	sink0_endofpacket;
output 	nxt_out_eop;
input 	cp_ready;
output 	in_data_reg_60;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_6;
input 	write_cp_data_69;
input 	write_cp_data_68;
input 	write_cp_data_67;
input 	write_cp_data_66;
input 	write_cp_data_65;
input 	WideNor0;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	base_address_3;
input 	base_address_2;
input 	out_data_1;
input 	out_data_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~2_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~2_combout ;
wire \Selector1~0_combout ;
wire \Selector1~3_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~7_combout ;
wire \d0_int_bytes_remaining[2]~8_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~5_combout ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~1_combout ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~5_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~6_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \d0_int_nxt_addr[3]~1_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~2_combout ;
wire \d0_int_nxt_addr[2]~3_combout ;
wire \in_eop_reg~q ;


terminal_qsys_altera_merlin_address_alignment_1 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_77(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold1),
	.datac(!out_valid_reg1),
	.datad(!write),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "on";
defparam \nxt_in_ready~1 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_ready_hold(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_hold1),
	.prn(vcc));
defparam in_ready_hold.is_wysiwyg = "true";
defparam in_ready_hold.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[59] (
	.clk(clk_clk),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!write),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(clk_clk),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(clk_clk),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(clk_clk),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(clk_clk),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(clk_clk),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(clk_clk),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(clk_clk),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(clk_clk),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(clk_clk),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(clk_clk),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(clk_clk),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(clk_clk),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(clk_clk),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(clk_clk),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(clk_clk),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(clk_clk),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(clk_clk),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(clk_clk),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(clk_clk),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(clk_clk),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(clk_clk),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(clk_clk),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(clk_clk),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(clk_clk),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(clk_clk),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!write),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[60] (
	.clk(clk_clk),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(clk_clk),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(clk_clk),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(clk_clk),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(clk_clk),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(clk_clk),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(clk_clk),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[100] (
	.clk(clk_clk),
	.d(sink0_data[100]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_100),
	.prn(vcc));
defparam \in_data_reg[100] .is_wysiwyg = "true";
defparam \in_data_reg[100] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(clk_clk),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(clk_clk),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(clk_clk),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold1),
	.datab(!sink0_data[59]),
	.datac(!Equal3),
	.datad(!Equal4),
	.datae(!src3_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold1),
	.datab(!sink0_data[59]),
	.datac(!Equal3),
	.datad(!Equal4),
	.datae(!src3_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[4]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[3]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[5]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!\WideOr0~combout ),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[60]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BF370A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h4454445444544454;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!sink0_data[60]),
	.datab(!\in_valid~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h1111111111111111;
defparam \Selector1~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~7 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~7 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~8 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~5 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~5 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[59]),
	.datad(!Add2),
	.datae(!write_cp_data_67),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'hCCDDCFDF00110313;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!Add21),
	.datad(!write_cp_data_68),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h0537053705370537;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!Add22),
	.datad(!write_cp_data_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h0537053705370537;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[4]~4_combout ),
	.datab(!\d0_int_bytes_remaining[3]~6_combout ),
	.datac(!\d0_int_bytes_remaining[2]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0808080808080808;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~2_combout ),
	.datab(!\Selector1~0_combout ),
	.datac(!\Selector1~3_combout ),
	.datad(!\d0_int_bytes_remaining[6]~1_combout ),
	.datae(!\d0_int_bytes_remaining[5]~3_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hA2A2A2A2FFA2A2A2;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[60]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[59]),
	.datae(!\in_valid~combout ),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h3030777530303330;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!\in_valid~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0707070707070707;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\Selector3~0_combout ),
	.datab(!\WideOr0~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h1111111111111111;
defparam \Selector3~1 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[71]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~5 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~5 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~5 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[0]~q ),
	.datac(!\d0_int_nxt_addr[0]~6_combout ),
	.datad(!sink0_data[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0D080D080D080D08;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~5_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~6 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~6 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!\ShiftLeft0~3_combout ),
	.datab(!\d0_int_nxt_addr[1]~4_combout ),
	.datac(!\int_nxt_addr_reg[1]~q ),
	.datad(!\in_burstwrap_reg[1]~q ),
	.datae(!\Add0~9_sumout ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h0F0F0FFF11111111;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[73]),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\int_nxt_addr_reg[3]~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~1 .lut_mask = 64'h0022AAAA5577FFFF;
defparam \d0_int_nxt_addr[3]~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[72]),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~2 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~2 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~5_sumout ),
	.datac(gnd),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\int_nxt_addr_reg[2]~q ),
	.dataf(!\d0_int_nxt_addr[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~3 .lut_mask = 64'h0022AAAA5577FFFF;
defparam \d0_int_nxt_addr[2]~3 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module terminal_qsys_altera_merlin_address_alignment_1 (
	new_burst_reg,
	src_data_77,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_77;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_77),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_adapter_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	nxt_in_ready,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	out_valid_reg,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_59,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sop_enable,
	Equal3,
	Equal31,
	saved_grant_0,
	in_data_reg_0,
	altera_reset_synchronizer_int_chain_out,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	Add2,
	Add21,
	Add22,
	burst_bytecount_6,
	write_cp_data_69,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_2,
	write_cp_data_65,
	WideNor0,
	src2_valid,
	src_valid,
	src_payload_0,
	nxt_out_eop,
	cp_ready,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	base_address_3,
	base_address_2,
	src_payload,
	src_data_73,
	src_data_72,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	src_data_77,
	out_data_1,
	src_data_71,
	out_data_0,
	src_data_70,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
output 	nxt_in_ready;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_59;
input 	write;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	sop_enable;
input 	Equal3;
input 	Equal31;
input 	saved_grant_0;
output 	in_data_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	Add2;
input 	Add21;
input 	Add22;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	burst_bytecount_4;
input 	write_cp_data_67;
input 	burst_bytecount_3;
input 	write_cp_data_66;
input 	burst_bytecount_2;
input 	write_cp_data_65;
output 	WideNor0;
input 	src2_valid;
input 	src_valid;
input 	src_payload_0;
output 	nxt_out_eop;
input 	cp_ready;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	base_address_3;
input 	base_address_2;
input 	src_payload;
input 	src_data_73;
input 	src_data_72;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_100;
input 	src_data_101;
input 	src_data_102;
input 	src_data_103;
input 	src_data_77;
input 	out_data_1;
input 	src_data_71;
input 	out_data_0;
input 	src_data_70;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_adapter_13_1_1 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_103,src_data_102,src_data_101,src_data_100,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,src_data_77,gnd,gnd,gnd,
src_data_73,src_data_72,src_data_71,src_data_70,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,src_payload31,src_payload30,src_payload29,
src_payload28,src_payload27,src_payload26,src_payload25,src_payload24,src_payload23,src_payload22,src_payload21,src_payload20,src_payload19,src_payload18,src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload11,src_payload10,
src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_59(in_data_reg_59),
	.write(write),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.sop_enable(sop_enable),
	.Equal3(Equal3),
	.Equal31(Equal31),
	.in_data_reg_0(in_data_reg_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.in_data_reg_10(in_data_reg_10),
	.in_data_reg_11(in_data_reg_11),
	.in_data_reg_12(in_data_reg_12),
	.in_data_reg_13(in_data_reg_13),
	.in_data_reg_14(in_data_reg_14),
	.in_data_reg_15(in_data_reg_15),
	.in_data_reg_16(in_data_reg_16),
	.in_data_reg_17(in_data_reg_17),
	.in_data_reg_18(in_data_reg_18),
	.in_data_reg_19(in_data_reg_19),
	.in_data_reg_20(in_data_reg_20),
	.in_data_reg_21(in_data_reg_21),
	.in_data_reg_22(in_data_reg_22),
	.in_data_reg_23(in_data_reg_23),
	.in_data_reg_24(in_data_reg_24),
	.in_data_reg_25(in_data_reg_25),
	.in_data_reg_26(in_data_reg_26),
	.in_data_reg_27(in_data_reg_27),
	.in_data_reg_28(in_data_reg_28),
	.in_data_reg_29(in_data_reg_29),
	.in_data_reg_30(in_data_reg_30),
	.in_data_reg_31(in_data_reg_31),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.burst_bytecount_6(burst_bytecount_6),
	.write_cp_data_69(write_cp_data_69),
	.burst_bytecount_5(burst_bytecount_5),
	.write_cp_data_68(write_cp_data_68),
	.burst_bytecount_4(burst_bytecount_4),
	.write_cp_data_67(write_cp_data_67),
	.burst_bytecount_3(burst_bytecount_3),
	.write_cp_data_66(write_cp_data_66),
	.burst_bytecount_2(burst_bytecount_2),
	.write_cp_data_65(write_cp_data_65),
	.WideNor0(WideNor0),
	.src2_valid(src2_valid),
	.src_valid(src_valid),
	.sink0_endofpacket(src_payload_0),
	.nxt_out_eop(nxt_out_eop),
	.cp_ready(cp_ready),
	.in_data_reg_60(in_data_reg_60),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_100(in_data_reg_100),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.base_address_3(base_address_3),
	.base_address_2(base_address_2),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_merlin_burst_adapter_13_1_1 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	nxt_in_ready,
	in_ready_hold,
	sink0_data,
	stateST_COMP_TRANS,
	out_valid_reg1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_59,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	sop_enable,
	Equal3,
	Equal31,
	in_data_reg_0,
	altera_reset_synchronizer_int_chain_out,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	in_data_reg_10,
	in_data_reg_11,
	in_data_reg_12,
	in_data_reg_13,
	in_data_reg_14,
	in_data_reg_15,
	in_data_reg_16,
	in_data_reg_17,
	in_data_reg_18,
	in_data_reg_19,
	in_data_reg_20,
	in_data_reg_21,
	in_data_reg_22,
	in_data_reg_23,
	in_data_reg_24,
	in_data_reg_25,
	in_data_reg_26,
	in_data_reg_27,
	in_data_reg_28,
	in_data_reg_29,
	in_data_reg_30,
	in_data_reg_31,
	Add2,
	Add21,
	Add22,
	burst_bytecount_6,
	write_cp_data_69,
	burst_bytecount_5,
	write_cp_data_68,
	burst_bytecount_4,
	write_cp_data_67,
	burst_bytecount_3,
	write_cp_data_66,
	burst_bytecount_2,
	write_cp_data_65,
	WideNor0,
	src2_valid,
	src_valid,
	sink0_endofpacket,
	nxt_out_eop,
	cp_ready,
	in_data_reg_60,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	base_address_3,
	base_address_2,
	out_data_1,
	out_data_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
output 	nxt_in_ready;
input 	in_ready_hold;
input 	[115:0] sink0_data;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_59;
input 	write;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	sop_enable;
input 	Equal3;
input 	Equal31;
output 	in_data_reg_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
output 	in_data_reg_10;
output 	in_data_reg_11;
output 	in_data_reg_12;
output 	in_data_reg_13;
output 	in_data_reg_14;
output 	in_data_reg_15;
output 	in_data_reg_16;
output 	in_data_reg_17;
output 	in_data_reg_18;
output 	in_data_reg_19;
output 	in_data_reg_20;
output 	in_data_reg_21;
output 	in_data_reg_22;
output 	in_data_reg_23;
output 	in_data_reg_24;
output 	in_data_reg_25;
output 	in_data_reg_26;
output 	in_data_reg_27;
output 	in_data_reg_28;
output 	in_data_reg_29;
output 	in_data_reg_30;
output 	in_data_reg_31;
input 	Add2;
input 	Add21;
input 	Add22;
input 	burst_bytecount_6;
input 	write_cp_data_69;
input 	burst_bytecount_5;
input 	write_cp_data_68;
input 	burst_bytecount_4;
input 	write_cp_data_67;
input 	burst_bytecount_3;
input 	write_cp_data_66;
input 	burst_bytecount_2;
input 	write_cp_data_65;
output 	WideNor0;
input 	src2_valid;
input 	src_valid;
input 	sink0_endofpacket;
output 	nxt_out_eop;
input 	cp_ready;
output 	in_data_reg_60;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	base_address_3;
input 	base_address_2;
input 	out_data_1;
input 	out_data_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \in_valid~combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~1_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~5_combout ;
wire \WideOr0~combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \nxt_in_ready~0_combout ;
wire \Selector1~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~7_combout ;
wire \d0_int_bytes_remaining[2]~8_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~5_combout ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~2_combout ;
wire \WideNor0~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~5_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~6_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \d0_int_nxt_addr[3]~1_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~2_combout ;
wire \d0_int_nxt_addr[2]~3_combout ;
wire \in_eop_reg~q ;


terminal_qsys_altera_merlin_address_alignment_2 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_77(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!write),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "on";
defparam \nxt_in_ready~2 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~2 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[59] (
	.clk(clk_clk),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!write),
	.datad(!\nxt_in_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h8A008A008A008A00;
defparam \nxt_in_ready~1 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(clk_clk),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(clk_clk),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(clk_clk),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

dffeas \in_data_reg[10] (
	.clk(clk_clk),
	.d(sink0_data[10]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_10),
	.prn(vcc));
defparam \in_data_reg[10] .is_wysiwyg = "true";
defparam \in_data_reg[10] .power_up = "low";

dffeas \in_data_reg[11] (
	.clk(clk_clk),
	.d(sink0_data[11]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_11),
	.prn(vcc));
defparam \in_data_reg[11] .is_wysiwyg = "true";
defparam \in_data_reg[11] .power_up = "low";

dffeas \in_data_reg[12] (
	.clk(clk_clk),
	.d(sink0_data[12]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_12),
	.prn(vcc));
defparam \in_data_reg[12] .is_wysiwyg = "true";
defparam \in_data_reg[12] .power_up = "low";

dffeas \in_data_reg[13] (
	.clk(clk_clk),
	.d(sink0_data[13]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_13),
	.prn(vcc));
defparam \in_data_reg[13] .is_wysiwyg = "true";
defparam \in_data_reg[13] .power_up = "low";

dffeas \in_data_reg[14] (
	.clk(clk_clk),
	.d(sink0_data[14]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_14),
	.prn(vcc));
defparam \in_data_reg[14] .is_wysiwyg = "true";
defparam \in_data_reg[14] .power_up = "low";

dffeas \in_data_reg[15] (
	.clk(clk_clk),
	.d(sink0_data[15]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_15),
	.prn(vcc));
defparam \in_data_reg[15] .is_wysiwyg = "true";
defparam \in_data_reg[15] .power_up = "low";

dffeas \in_data_reg[16] (
	.clk(clk_clk),
	.d(sink0_data[16]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_16),
	.prn(vcc));
defparam \in_data_reg[16] .is_wysiwyg = "true";
defparam \in_data_reg[16] .power_up = "low";

dffeas \in_data_reg[17] (
	.clk(clk_clk),
	.d(sink0_data[17]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_17),
	.prn(vcc));
defparam \in_data_reg[17] .is_wysiwyg = "true";
defparam \in_data_reg[17] .power_up = "low";

dffeas \in_data_reg[18] (
	.clk(clk_clk),
	.d(sink0_data[18]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_18),
	.prn(vcc));
defparam \in_data_reg[18] .is_wysiwyg = "true";
defparam \in_data_reg[18] .power_up = "low";

dffeas \in_data_reg[19] (
	.clk(clk_clk),
	.d(sink0_data[19]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_19),
	.prn(vcc));
defparam \in_data_reg[19] .is_wysiwyg = "true";
defparam \in_data_reg[19] .power_up = "low";

dffeas \in_data_reg[20] (
	.clk(clk_clk),
	.d(sink0_data[20]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_20),
	.prn(vcc));
defparam \in_data_reg[20] .is_wysiwyg = "true";
defparam \in_data_reg[20] .power_up = "low";

dffeas \in_data_reg[21] (
	.clk(clk_clk),
	.d(sink0_data[21]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_21),
	.prn(vcc));
defparam \in_data_reg[21] .is_wysiwyg = "true";
defparam \in_data_reg[21] .power_up = "low";

dffeas \in_data_reg[22] (
	.clk(clk_clk),
	.d(sink0_data[22]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_22),
	.prn(vcc));
defparam \in_data_reg[22] .is_wysiwyg = "true";
defparam \in_data_reg[22] .power_up = "low";

dffeas \in_data_reg[23] (
	.clk(clk_clk),
	.d(sink0_data[23]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_23),
	.prn(vcc));
defparam \in_data_reg[23] .is_wysiwyg = "true";
defparam \in_data_reg[23] .power_up = "low";

dffeas \in_data_reg[24] (
	.clk(clk_clk),
	.d(sink0_data[24]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_24),
	.prn(vcc));
defparam \in_data_reg[24] .is_wysiwyg = "true";
defparam \in_data_reg[24] .power_up = "low";

dffeas \in_data_reg[25] (
	.clk(clk_clk),
	.d(sink0_data[25]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_25),
	.prn(vcc));
defparam \in_data_reg[25] .is_wysiwyg = "true";
defparam \in_data_reg[25] .power_up = "low";

dffeas \in_data_reg[26] (
	.clk(clk_clk),
	.d(sink0_data[26]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_26),
	.prn(vcc));
defparam \in_data_reg[26] .is_wysiwyg = "true";
defparam \in_data_reg[26] .power_up = "low";

dffeas \in_data_reg[27] (
	.clk(clk_clk),
	.d(sink0_data[27]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_27),
	.prn(vcc));
defparam \in_data_reg[27] .is_wysiwyg = "true";
defparam \in_data_reg[27] .power_up = "low";

dffeas \in_data_reg[28] (
	.clk(clk_clk),
	.d(sink0_data[28]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_28),
	.prn(vcc));
defparam \in_data_reg[28] .is_wysiwyg = "true";
defparam \in_data_reg[28] .power_up = "low";

dffeas \in_data_reg[29] (
	.clk(clk_clk),
	.d(sink0_data[29]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_29),
	.prn(vcc));
defparam \in_data_reg[29] .is_wysiwyg = "true";
defparam \in_data_reg[29] .power_up = "low";

dffeas \in_data_reg[30] (
	.clk(clk_clk),
	.d(sink0_data[30]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_30),
	.prn(vcc));
defparam \in_data_reg[30] .is_wysiwyg = "true";
defparam \in_data_reg[30] .power_up = "low";

dffeas \in_data_reg[31] (
	.clk(clk_clk),
	.d(sink0_data[31]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_31),
	.prn(vcc));
defparam \in_data_reg[31] .is_wysiwyg = "true";
defparam \in_data_reg[31] .power_up = "low";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sop_enable),
	.datab(!burst_bytecount_6),
	.datac(!burst_bytecount_5),
	.datad(!burst_bytecount_3),
	.datae(!burst_bytecount_2),
	.dataf(!burst_bytecount_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideNor0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h4000000000000000;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!write),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[60] (
	.clk(clk_clk),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(clk_clk),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(clk_clk),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(clk_clk),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(clk_clk),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(clk_clk),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(clk_clk),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[100] (
	.clk(clk_clk),
	.d(sink0_data[100]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_100),
	.prn(vcc));
defparam \in_data_reg[100] .is_wysiwyg = "true";
defparam \in_data_reg[100] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(clk_clk),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(clk_clk),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(clk_clk),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

cyclonev_lcell_comb in_valid(
	.dataa(!in_ready_hold),
	.datab(!sink0_data[59]),
	.datac(!Equal3),
	.datad(!Equal31),
	.datae(!src2_valid),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam in_valid.extended_lut = "off";
defparam in_valid.lut_mask = 64'h0000000155555555;
defparam in_valid.shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[60]),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h005FCCFF005FCCFF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[59]),
	.datac(!Equal3),
	.datad(!Equal31),
	.datae(!src2_valid),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0000000100000000;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[2]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[6]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~1_combout ),
	.datac(!\in_valid~combout ),
	.datad(!\WideOr0~combout ),
	.datae(!\state.ST_UNCOMP_TRANS~q ),
	.dataf(!sink0_data[60]),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "on";
defparam \Selector2~2 .lut_mask = 64'h3B33BF370A00AA00;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!sink0_data[59]),
	.datad(!\in_valid~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h4454445444544454;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_in_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!sink0_data[60]),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!\nxt_in_ready~0_combout ),
	.datae(!\in_valid~combout ),
	.dataf(!\state.ST_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h0000555500001511;
defparam \Selector1~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~7 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~7 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~8 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~5 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~5 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[59]),
	.datad(!Add2),
	.datae(!\Add1~1_combout ),
	.dataf(!write_cp_data_67),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'hCCDD0011CFDF0313;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!Add21),
	.datad(!write_cp_data_68),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h0537053705370537;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!Add22),
	.datad(!write_cp_data_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h0537053705370537;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[3]~6_combout ),
	.datab(!\d0_int_bytes_remaining[2]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h2222222222222222;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\Selector1~1_combout ),
	.datac(!\d0_int_bytes_remaining[6]~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~3_combout ),
	.datae(!\d0_int_bytes_remaining[4]~4_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'h88888888F8888888;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!\state.ST_IDLE~q ),
	.datab(!\in_valid~combout ),
	.datac(!sink0_data[59]),
	.datad(!nxt_out_eop),
	.datae(!stateST_COMP_TRANS),
	.dataf(!sink0_data[60]),
	.datag(!\nxt_in_ready~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "on";
defparam \Selector1~2 .lut_mask = 64'h0000FF302232FF33;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~1 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~1 .extended_lut = "off";
defparam \WideNor0~1 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!\in_valid~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0707070707070707;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!\in_valid~combout ),
	.datae(!cp_ready),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h50FF44FF50FF44FF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\nxt_in_ready~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8888888888888888;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\Selector3~0_combout ),
	.datab(!\WideOr0~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h1111111111111111;
defparam \Selector3~1 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h10BA101010BA1010;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[1]~q ),
	.datae(!\in_size_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[71]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~5 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~5 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~5 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[0]~q ),
	.datac(!\d0_int_nxt_addr[0]~6_combout ),
	.datad(!sink0_data[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0D080D080D080D08;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~5_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~6 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~6 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!\ShiftLeft0~3_combout ),
	.datab(!\d0_int_nxt_addr[1]~4_combout ),
	.datac(!\int_nxt_addr_reg[1]~q ),
	.datad(!\in_burstwrap_reg[1]~q ),
	.datae(!\Add0~9_sumout ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h0F0F0FFF11111111;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[73]),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\int_nxt_addr_reg[3]~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~1 .lut_mask = 64'h0022AAAA5577FFFF;
defparam \d0_int_nxt_addr[3]~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[72]),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~2 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~2 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~5_sumout ),
	.datac(gnd),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\int_nxt_addr_reg[2]~q ),
	.dataf(!\d0_int_nxt_addr[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~3 .lut_mask = 64'h0022AAAA5577FFFF;
defparam \d0_int_nxt_addr[2]~3 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module terminal_qsys_altera_merlin_address_alignment_2 (
	new_burst_reg,
	src_data_77,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_77;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_77),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_adapter_2 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	nxt_in_ready,
	in_ready_hold,
	saved_grant_1,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_59,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	Add2,
	Add21,
	Add22,
	write_cp_data_69,
	write_cp_data_68,
	write_cp_data_67,
	write_cp_data_66,
	write_cp_data_65,
	WideNor0,
	src_valid,
	src_valid1,
	src_payload_0,
	nxt_out_eop,
	cp_ready,
	cp_ready1,
	in_data_reg_60,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	base_address_3,
	base_address_2,
	src_payload,
	src_data_73,
	src_data_72,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	nxt_in_ready2,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	src_data_77,
	out_data_1,
	src_data_71,
	out_data_0,
	src_data_70,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
output 	nxt_in_ready;
input 	in_ready_hold;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
output 	out_valid_reg;
input 	mem_used_1;
output 	in_narrow_reg;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_59;
input 	write;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
input 	Add2;
input 	Add21;
input 	Add22;
input 	write_cp_data_69;
input 	write_cp_data_68;
input 	write_cp_data_67;
input 	write_cp_data_66;
input 	write_cp_data_65;
input 	WideNor0;
input 	src_valid;
input 	src_valid1;
input 	src_payload_0;
output 	nxt_out_eop;
input 	cp_ready;
input 	cp_ready1;
output 	in_data_reg_60;
input 	src_data_78;
input 	src_data_79;
input 	src_data_35;
input 	src_data_34;
input 	src_data_33;
input 	src_data_32;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	base_address_3;
input 	base_address_2;
input 	src_payload;
input 	src_data_73;
input 	src_data_72;
input 	src_payload1;
input 	src_payload2;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
output 	nxt_in_ready2;
input 	src_data_92;
input 	src_data_93;
input 	src_data_94;
input 	src_data_95;
input 	src_data_96;
input 	src_data_97;
input 	src_data_98;
input 	src_data_99;
input 	src_data_100;
input 	src_data_101;
input 	src_data_102;
input 	src_data_103;
input 	src_data_77;
input 	out_data_1;
input 	src_data_71;
input 	out_data_0;
input 	src_data_70;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_adapter_13_1_2 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.nxt_in_ready(nxt_in_ready),
	.in_ready_hold(in_ready_hold),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_103,src_data_102,src_data_101,src_data_100,src_data_99,src_data_98,src_data_97,src_data_96,src_data_95,src_data_94,src_data_93,src_data_92,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_79,src_data_78,src_data_77,gnd,gnd,gnd,
src_data_73,src_data_72,src_data_71,src_data_70,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,saved_grant_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_35,src_data_34,src_data_33,src_data_32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload9,src_payload8,src_payload7,src_payload6,src_payload5,src_payload4,src_payload3,src_payload2,src_payload1,src_payload}),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.out_valid_reg1(out_valid_reg),
	.mem_used_1(mem_used_1),
	.in_narrow_reg1(in_narrow_reg),
	.in_byteen_reg_3(in_byteen_reg_3),
	.in_byteen_reg_2(in_byteen_reg_2),
	.in_byteen_reg_1(in_byteen_reg_1),
	.in_byteen_reg_0(in_byteen_reg_0),
	.in_data_reg_59(in_data_reg_59),
	.write(write),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.in_data_reg_0(in_data_reg_0),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_1(in_data_reg_1),
	.in_data_reg_2(in_data_reg_2),
	.in_data_reg_3(in_data_reg_3),
	.in_data_reg_4(in_data_reg_4),
	.in_data_reg_5(in_data_reg_5),
	.in_data_reg_6(in_data_reg_6),
	.in_data_reg_7(in_data_reg_7),
	.in_data_reg_8(in_data_reg_8),
	.in_data_reg_9(in_data_reg_9),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.write_cp_data_69(write_cp_data_69),
	.write_cp_data_68(write_cp_data_68),
	.write_cp_data_67(write_cp_data_67),
	.write_cp_data_66(write_cp_data_66),
	.write_cp_data_65(write_cp_data_65),
	.WideNor0(WideNor0),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.sink0_endofpacket(src_payload_0),
	.nxt_out_eop(nxt_out_eop),
	.cp_ready(cp_ready),
	.cp_ready1(cp_ready1),
	.in_data_reg_60(in_data_reg_60),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_100(in_data_reg_100),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.base_address_3(base_address_3),
	.base_address_2(base_address_2),
	.nxt_in_ready2(nxt_in_ready2),
	.out_data_1(out_data_1),
	.out_data_0(out_data_0),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_merlin_burst_adapter_13_1_2 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	nxt_in_ready,
	in_ready_hold,
	sink0_data,
	stateST_COMP_TRANS,
	out_valid_reg1,
	mem_used_1,
	in_narrow_reg1,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	in_data_reg_59,
	write,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	altera_reset_synchronizer_int_chain_out,
	in_data_reg_0,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	in_data_reg_1,
	in_data_reg_2,
	in_data_reg_3,
	in_data_reg_4,
	in_data_reg_5,
	in_data_reg_6,
	in_data_reg_7,
	in_data_reg_8,
	in_data_reg_9,
	Add2,
	Add21,
	Add22,
	write_cp_data_69,
	write_cp_data_68,
	write_cp_data_67,
	write_cp_data_66,
	write_cp_data_65,
	WideNor0,
	src_valid,
	src_valid1,
	sink0_endofpacket,
	nxt_out_eop,
	cp_ready,
	cp_ready1,
	in_data_reg_60,
	out_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	base_address_3,
	base_address_2,
	nxt_in_ready2,
	out_data_1,
	out_data_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
output 	nxt_in_ready;
input 	in_ready_hold;
input 	[115:0] sink0_data;
output 	stateST_COMP_TRANS;
output 	out_valid_reg1;
input 	mem_used_1;
output 	in_narrow_reg1;
output 	in_byteen_reg_3;
output 	in_byteen_reg_2;
output 	in_byteen_reg_1;
output 	in_byteen_reg_0;
output 	in_data_reg_59;
input 	write;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	altera_reset_synchronizer_int_chain_out;
output 	in_data_reg_0;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_1;
output 	in_data_reg_2;
output 	in_data_reg_3;
output 	in_data_reg_4;
output 	in_data_reg_5;
output 	in_data_reg_6;
output 	in_data_reg_7;
output 	in_data_reg_8;
output 	in_data_reg_9;
input 	Add2;
input 	Add21;
input 	Add22;
input 	write_cp_data_69;
input 	write_cp_data_68;
input 	write_cp_data_67;
input 	write_cp_data_66;
input 	write_cp_data_65;
input 	WideNor0;
input 	src_valid;
input 	src_valid1;
input 	sink0_endofpacket;
output 	nxt_out_eop;
input 	cp_ready;
input 	cp_ready1;
output 	in_data_reg_60;
output 	out_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	base_address_3;
input 	base_address_2;
output 	nxt_in_ready2;
input 	out_data_1;
input 	out_data_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \Selector3~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideOr0~0_combout ;
wire \Selector0~0_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_IDLE~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[2]~7_combout ;
wire \d0_int_bytes_remaining[2]~8_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~5_combout ;
wire \d0_int_bytes_remaining[3]~6_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~4_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \d0_int_bytes_remaining[5]~3_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~0_combout ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \Equal0~0_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \Selector1~3_combout ;
wire \WideNor0~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \LessThan0~0_combout ;
wire \Selector3~1_combout ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \ShiftLeft0~3_combout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~4_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \d0_int_nxt_addr[0]~5_combout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~6_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~7_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \d0_int_nxt_addr[3]~1_combout ;
wire \Add0~5_sumout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \d0_int_nxt_addr[2]~2_combout ;
wire \d0_int_nxt_addr[2]~3_combout ;
wire \in_eop_reg~q ;


terminal_qsys_altera_merlin_address_alignment_3 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_data_77(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.ShiftLeft0(\ShiftLeft0~3_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

cyclonev_lcell_comb \nxt_in_ready~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!in_ready_hold),
	.datac(!out_valid_reg1),
	.datad(!write),
	.datae(!stateST_COMP_TRANS),
	.dataf(!\new_burst_reg~q ),
	.datag(!stateST_UNCOMP_WR_SUBBURST),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~2 .extended_lut = "on";
defparam \nxt_in_ready~2 .lut_mask = 64'h2020F0F02020F0FF;
defparam \nxt_in_ready~2 .shared_arith = "off";

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

dffeas \in_byteen_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[35]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_3),
	.prn(vcc));
defparam \in_byteen_reg[3] .is_wysiwyg = "true";
defparam \in_byteen_reg[3] .power_up = "low";

dffeas \in_byteen_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[34]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_2),
	.prn(vcc));
defparam \in_byteen_reg[2] .is_wysiwyg = "true";
defparam \in_byteen_reg[2] .power_up = "low";

dffeas \in_byteen_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[33]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_1),
	.prn(vcc));
defparam \in_byteen_reg[1] .is_wysiwyg = "true";
defparam \in_byteen_reg[1] .power_up = "low";

dffeas \in_byteen_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[32]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_byteen_reg_0),
	.prn(vcc));
defparam \in_byteen_reg[0] .is_wysiwyg = "true";
defparam \in_byteen_reg[0] .power_up = "low";

dffeas \in_data_reg[59] (
	.clk(clk_clk),
	.d(sink0_data[59]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_59),
	.prn(vcc));
defparam \in_data_reg[59] .is_wysiwyg = "true";
defparam \in_data_reg[59] .power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!out_valid_reg1),
	.datac(!write),
	.datad(!\state.ST_UNCOMP_TRANS~q ),
	.datae(!stateST_UNCOMP_WR_SUBBURST),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h008A8A8A008A8A8A;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas \in_data_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_0),
	.prn(vcc));
defparam \in_data_reg[0] .is_wysiwyg = "true";
defparam \in_data_reg[0] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_1),
	.prn(vcc));
defparam \in_data_reg[1] .is_wysiwyg = "true";
defparam \in_data_reg[1] .power_up = "low";

dffeas \in_data_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_2),
	.prn(vcc));
defparam \in_data_reg[2] .is_wysiwyg = "true";
defparam \in_data_reg[2] .power_up = "low";

dffeas \in_data_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_3),
	.prn(vcc));
defparam \in_data_reg[3] .is_wysiwyg = "true";
defparam \in_data_reg[3] .power_up = "low";

dffeas \in_data_reg[4] (
	.clk(clk_clk),
	.d(sink0_data[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_4),
	.prn(vcc));
defparam \in_data_reg[4] .is_wysiwyg = "true";
defparam \in_data_reg[4] .power_up = "low";

dffeas \in_data_reg[5] (
	.clk(clk_clk),
	.d(sink0_data[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_5),
	.prn(vcc));
defparam \in_data_reg[5] .is_wysiwyg = "true";
defparam \in_data_reg[5] .power_up = "low";

dffeas \in_data_reg[6] (
	.clk(clk_clk),
	.d(sink0_data[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_6),
	.prn(vcc));
defparam \in_data_reg[6] .is_wysiwyg = "true";
defparam \in_data_reg[6] .power_up = "low";

dffeas \in_data_reg[7] (
	.clk(clk_clk),
	.d(sink0_data[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_7),
	.prn(vcc));
defparam \in_data_reg[7] .is_wysiwyg = "true";
defparam \in_data_reg[7] .power_up = "low";

dffeas \in_data_reg[8] (
	.clk(clk_clk),
	.d(sink0_data[8]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_8),
	.prn(vcc));
defparam \in_data_reg[8] .is_wysiwyg = "true";
defparam \in_data_reg[8] .power_up = "low";

dffeas \in_data_reg[9] (
	.clk(clk_clk),
	.d(sink0_data[9]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_9),
	.prn(vcc));
defparam \in_data_reg[9] .is_wysiwyg = "true";
defparam \in_data_reg[9] .power_up = "low";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!\in_eop_reg~q ),
	.datab(!stateST_COMP_TRANS),
	.datac(!\new_burst_reg~q ),
	.datad(!write),
	.datae(!\in_bytecount_reg_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h4447774744477747;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \in_data_reg[60] (
	.clk(clk_clk),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(clk_clk),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(clk_clk),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(clk_clk),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(clk_clk),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(clk_clk),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(clk_clk),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[100] (
	.clk(clk_clk),
	.d(sink0_data[100]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_100),
	.prn(vcc));
defparam \in_data_reg[100] .is_wysiwyg = "true";
defparam \in_data_reg[100] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(clk_clk),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(clk_clk),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(clk_clk),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h8888888888888888;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!out_valid_reg1),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h1111111111111111;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_3),
	.datab(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datac(!out_uncomp_byte_cnt_reg_2),
	.datad(!out_uncomp_byte_cnt_reg_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h2000200020002000;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h04FEAE5404FEAE54;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_UNCOMP_TRANS~q ),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .lut_mask = 64'h0404AE04FEFE54FE;
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(!out_uncomp_byte_cnt_reg_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .lut_mask = 64'h00E40044FF4EFFEE;
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h8080808080808080;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!sink0_data[59]),
	.datab(!src_valid1),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!\state.ST_IDLE~q ),
	.dataf(!in_ready_hold),
	.datag(!sink0_data[60]),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "on";
defparam \Selector0~0 .lut_mask = 64'h0000F0F0135FF3FF;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!out_valid_reg1),
	.datab(!write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!stateST_UNCOMP_WR_SUBBURST),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0001555500010101;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!sink0_data[60]),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datac(!\Selector3~0_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.datae(!\WideOr0~0_combout ),
	.dataf(!\Selector2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'h00000C00AAAAAEAA;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!nxt_out_eop),
	.datad(!sink0_data[59]),
	.datae(!src_valid),
	.dataf(!src_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h3030313031303130;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!nxt_out_eop),
	.datac(!\state.ST_UNCOMP_TRANS~q ),
	.datad(!stateST_UNCOMP_WR_SUBBURST),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h0000A8880000A888;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!in_ready_hold),
	.datab(!sink0_data[60]),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'h0111011101110111;
defparam \Selector1~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~7 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!write_cp_data_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~7 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~7 .lut_mask = 64'h2F222F222F222F22;
defparam \d0_int_bytes_remaining[2]~7 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~8 (
	.dataa(!\new_burst_reg~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\int_bytes_remaining_reg[2]~q ),
	.datad(!\d0_int_bytes_remaining[2]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~8 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~8 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[2]~8 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~5 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!sink0_data[60]),
	.datad(!sink0_data[59]),
	.datae(!write_cp_data_66),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~5 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~5 .lut_mask = 64'h060606FF060606FF;
defparam \d0_int_bytes_remaining[3]~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(!\d0_int_bytes_remaining[3]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~6 .extended_lut = "off";
defparam \d0_int_bytes_remaining[3]~6 .lut_mask = 64'h28227D7728227D77;
defparam \d0_int_bytes_remaining[3]~6 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~4 (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[59]),
	.datad(!Add2),
	.datae(!write_cp_data_67),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~4 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~4 .lut_mask = 64'hCCDDCFDF00110313;
defparam \d0_int_bytes_remaining[4]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h0800080008000800;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!Add21),
	.datad(!write_cp_data_68),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h0537053705370537;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[5]~q ),
	.datac(!\Add1~0_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~3 .lut_mask = 64'h287D287D287D287D;
defparam \d0_int_bytes_remaining[5]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!Add22),
	.datad(!write_cp_data_69),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~0 .lut_mask = 64'h0537053705370537;
defparam \d0_int_bytes_remaining[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\int_bytes_remaining_reg[6]~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!\d0_int_bytes_remaining[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h228277D7228277D7;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\d0_int_bytes_remaining[4]~4_combout ),
	.datab(!\d0_int_bytes_remaining[3]~6_combout ),
	.datac(!\d0_int_bytes_remaining[2]~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0808080808080808;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\Selector1~1_combout ),
	.datac(!\Selector1~2_combout ),
	.datad(!\d0_int_bytes_remaining[6]~1_combout ),
	.datae(!\d0_int_bytes_remaining[5]~3_combout ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hA2A2A2A2FFA2A2A2;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\Selector1~1_combout ),
	.datac(!\Selector1~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h5D5D5D5D5D5D5D5D;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \WideNor0~0 (
	.dataa(!sink0_data[60]),
	.datab(!sink0_data[59]),
	.datac(!WideNor0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor0~0 .extended_lut = "off";
defparam \WideNor0~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \WideNor0~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd (
	.dataa(!in_ready_hold),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready),
	.datad(!src_valid),
	.datae(!src_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd .lut_mask = 64'h0015151500151515;
defparam \NON_PIPELINED_INPUTS.load_next_cmd .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\WideNor0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!mem_used_1),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready),
	.datae(!cp_ready1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0B8B8B8F0B8B8B8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!\nxt_out_valid~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0555377705553777;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!sink0_data[78]),
	.datab(!sink0_data[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h8888888888888888;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\Selector3~0_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.datad(!\WideOr0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h3313331333133313;
defparam \Selector3~1 .shared_arith = "off";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h1010BA101010BA10;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[2]~q ),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'hEA404040EA404040;
defparam \ShiftLeft0~3 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!h2f_lw_ARADDR_1),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[71]),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~4 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~4 .extended_lut = "off";
defparam \ShiftLeft0~4 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~4 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~5 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!out_data_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~5 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~5 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[0]~5 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!\new_burst_reg~q ),
	.datab(!\in_burstwrap_reg[0]~q ),
	.datac(!\d0_int_nxt_addr[0]~6_combout ),
	.datad(!sink0_data[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0D080D080D080D08;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~6 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~13_sumout ),
	.datac(!\align_address_to_size|LessThan0~0_combout ),
	.datad(!\d0_int_nxt_addr[0]~5_combout ),
	.datae(!\int_nxt_addr_reg[0]~q ),
	.dataf(!\in_burstwrap_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~6 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~6 .lut_mask = 64'h0005AAAF2227AAAF;
defparam \d0_int_nxt_addr[0]~6 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~7 (
	.dataa(!\ShiftLeft0~3_combout ),
	.datab(!\d0_int_nxt_addr[1]~4_combout ),
	.datac(!\int_nxt_addr_reg[1]~q ),
	.datad(!\in_burstwrap_reg[1]~q ),
	.datae(!\Add0~9_sumout ),
	.dataf(!\new_burst_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~7 .extended_lut = "off";
defparam \d0_int_nxt_addr[1]~7 .lut_mask = 64'h0F0F0FFF11111111;
defparam \d0_int_nxt_addr[1]~7 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[73]),
	.datac(!\in_burstwrap_reg[3]~q ),
	.datad(!\d0_int_nxt_addr[3]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\int_nxt_addr_reg[3]~q ),
	.dataf(!\d0_int_nxt_addr[3]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~1 .lut_mask = 64'h0022AAAA5577FFFF;
defparam \d0_int_nxt_addr[3]~1 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[72]),
	.datac(!\in_burstwrap_reg[2]~q ),
	.datad(!\d0_int_nxt_addr[2]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h00E400E400E400E4;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~2 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!sink0_data[59]),
	.datad(!base_address_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~2 .lut_mask = 64'h111F111F111F111F;
defparam \d0_int_nxt_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!\Add0~5_sumout ),
	.datac(gnd),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\int_nxt_addr_reg[2]~q ),
	.dataf(!\d0_int_nxt_addr[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~3 .lut_mask = 64'h0022AAAA5577FFFF;
defparam \d0_int_nxt_addr[2]~3 .shared_arith = "off";

dffeas in_eop_reg(
	.clk(clk_clk),
	.d(sink0_endofpacket),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~combout ),
	.q(\in_eop_reg~q ),
	.prn(vcc));
defparam in_eop_reg.is_wysiwyg = "true";
defparam in_eop_reg.power_up = "low";

endmodule

module terminal_qsys_altera_merlin_address_alignment_3 (
	new_burst_reg,
	src_data_77,
	in_size_reg_0,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_data_77;
input 	in_size_reg_0;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_data_77),
	.datac(!in_size_reg_0),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_adapter_3 (
	h2f_lw_ARVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	in_ready_hold,
	has_pending_responses,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_60,
	in_narrow_reg,
	cp_ready,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	nxt_out_eop,
	Equal1,
	last_channel_0,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	int_nxt_addr_reg_dly_2,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	Selector11,
	src_payload,
	src_payload1,
	src_payload2,
	Selector12,
	nxt_out_burstwrap_1,
	nxt_out_burstwrap_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	in_ready_hold;
input 	has_pending_responses;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_60;
output 	in_narrow_reg;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
output 	nxt_out_eop;
input 	Equal1;
input 	last_channel_0;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	Selector11;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	Selector12;
input 	nxt_out_burstwrap_1;
input 	nxt_out_burstwrap_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_adapter_13_1_3 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARVALID_0(h2f_lw_ARVALID_0),
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload,
src_payload2,gnd,gnd,gnd,gnd,Selector11,Selector12,nxt_out_burstwrap_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.in_ready_hold(in_ready_hold),
	.has_pending_responses(has_pending_responses),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_60(in_data_reg_60),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.saved_grant_1(saved_grant_1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.nxt_out_eop(nxt_out_eop),
	.Equal1(Equal1),
	.last_channel_0(last_channel_0),
	.src_valid(src_valid),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready1(cp_ready1),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_100(in_data_reg_100),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_merlin_burst_adapter_13_1_3 (
	h2f_lw_ARVALID_0,
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	sink0_data,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	in_ready_hold,
	has_pending_responses,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_60,
	in_narrow_reg1,
	cp_ready,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	nxt_out_eop,
	Equal1,
	last_channel_0,
	src_valid,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_6,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	int_nxt_addr_reg_dly_2,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	nxt_out_burstwrap_1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	[115:0] sink0_data;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	in_ready_hold;
input 	has_pending_responses;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_60;
output 	in_narrow_reg1;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
output 	nxt_out_eop;
input 	Equal1;
input 	last_channel_0;
input 	src_valid;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_6;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	int_nxt_addr_reg_dly_2;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	nxt_out_burstwrap_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~1_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[2]~0_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[3]~4_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[4]~3_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \d0_int_bytes_remaining[6]~1_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[0]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~9_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~1_combout ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[1]~3_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[2]~0_combout ;


terminal_qsys_altera_merlin_address_alignment_4 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[78]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.ShiftLeft0(\ShiftLeft0~0_combout ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[60] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(!cp_ready),
	.datae(!\new_burst_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000004400000044;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!in_ready_hold),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h0000FF77A0A0F5F5;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!in_data_reg_60),
	.datad(!cp_ready),
	.datae(!\new_burst_reg~q ),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h0A0A0A4E5F1B5F5F;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(clk_clk),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(clk_clk),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(clk_clk),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(clk_clk),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(clk_clk),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(clk_clk),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[100] (
	.clk(clk_clk),
	.d(sink0_data[100]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_100),
	.prn(vcc));
defparam \in_data_reg[100] .is_wysiwyg = "true";
defparam \in_data_reg[100] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(clk_clk),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(clk_clk),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(clk_clk),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h0202020202020202;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_6),
	.datad(!out_uncomp_byte_cnt_reg_5),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!\Add4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .lut_mask = 64'h0F0F4E4EA50FE44E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[6]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[5]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[4]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[3]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!saved_grant_1),
	.datac(!in_ready_hold),
	.datad(!has_pending_responses),
	.datae(!Equal1),
	.dataf(!last_channel_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0000010000000101;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!nxt_out_eop),
	.datab(!\state.ST_IDLE~q ),
	.datac(!\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_data_reg_60),
	.datac(!nxt_out_eop),
	.datad(!\Selector2~0_combout ),
	.datae(!\state.ST_IDLE~q ),
	.dataf(!\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h50505050FFFF7755;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~1 (
	.dataa(!saved_grant_1),
	.datab(!in_ready_hold),
	.datac(!Equal1),
	.datad(!nxt_in_ready),
	.datae(!nxt_in_ready1),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~1 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~1 .lut_mask = 64'h0000000001010001;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~0 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~4 (
	.dataa(!\int_bytes_remaining_reg[2]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!saved_grant_1),
	.datad(!h2f_lw_ARLEN_1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_lw_ARLEN_0),
	.datag(!\int_bytes_remaining_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~4 .extended_lut = "on";
defparam \d0_int_bytes_remaining[3]~4 .lut_mask = 64'h2D2D000F2D2D0F00;
defparam \d0_int_bytes_remaining[3]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hB4F0B4F0B4F0B4F0;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~3 (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\Add1~1_combout ),
	.datad(!Add2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~3 .lut_mask = 64'hC0D1C0D1C0D1C0D1;
defparam \d0_int_bytes_remaining[4]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h4000400040004000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\int_bytes_remaining_reg[5]~q ),
	.datad(!\Add1~0_combout ),
	.datae(!Add21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h0CC01DD10CC01DD1;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~1 (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\int_bytes_remaining_reg[6]~q ),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~0_combout ),
	.dataf(!Add22),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~1 .lut_mask = 64'h0C0CC00C1D1DD11D;
defparam \d0_int_bytes_remaining[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\d0_int_bytes_remaining[2]~0_combout ),
	.datac(!\d0_int_bytes_remaining[6]~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(!\d0_int_bytes_remaining[4]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hBAAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!saved_grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\in_bytecount_reg_zero~q ),
	.datae(!\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.dataf(!cp_ready1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'h5500FFFF5140FFFF;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[72]),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\d0_int_nxt_addr[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[79]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[77]),
	.datae(!\in_size_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[78]),
	.datac(!\in_size_reg[1]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~3_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\in_size_reg[1]~q ),
	.datab(!sink0_data[78]),
	.datac(!sink0_data[79]),
	.datad(!\in_size_reg[0]~q ),
	.datae(!\new_burst_reg~q ),
	.dataf(!sink0_data[77]),
	.datag(!\in_size_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "on";
defparam \ShiftLeft0~2 .lut_mask = 64'h00A0000000A0C0C0;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~1_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(!\d0_int_nxt_addr[0]~2_combout ),
	.datae(!sink0_data[70]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h00F300E200F300E2;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~1 (
	.dataa(!\Add0~9_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~1 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(!\d0_int_nxt_addr[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~3 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~5_sumout ),
	.datac(!saved_grant_1),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_lw_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~3 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~3 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~0 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_address_alignment_4 (
	new_burst_reg,
	src_payload,
	in_size_reg_1,
	ShiftLeft0,
	LessThan0)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_1;
input 	ShiftLeft0;
output 	LessThan0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_1),
	.datad(!ShiftLeft0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_adapter_4 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	in_ready_hold,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_60,
	in_narrow_reg,
	cp_ready,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	nxt_out_eop,
	Equal2,
	src_valid,
	src_valid1,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	Selector10,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Selector12,
	src_payload,
	src_payload1,
	src_payload2,
	nxt_out_burstwrap_1,
	nxt_out_burstwrap_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_60;
output 	in_narrow_reg;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
output 	nxt_out_eop;
input 	Equal2;
input 	src_valid;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	Selector10;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Selector12;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
input 	nxt_out_burstwrap_1;
input 	nxt_out_burstwrap_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_adapter_13_1_4 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload2,
src_payload,gnd,gnd,gnd,Selector10,Selector11,Selector12,nxt_out_burstwrap_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,saved_grant_1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.in_ready_hold(in_ready_hold),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_60(in_data_reg_60),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Decoder1(Decoder1),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.nxt_out_eop(nxt_out_eop),
	.Equal2(Equal2),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.cp_ready1(cp_ready1),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_100(in_data_reg_100),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_merlin_burst_adapter_13_1_4 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	sink0_data,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	in_ready_hold,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_60,
	in_narrow_reg1,
	cp_ready,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	altera_reset_synchronizer_int_chain_out,
	Decoder1,
	Add2,
	Add21,
	Add22,
	nxt_out_eop,
	Equal2,
	src_valid,
	src_valid1,
	out_byte_cnt_reg_2,
	cp_ready1,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	nxt_out_burstwrap_1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	[115:0] sink0_data;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	in_ready_hold;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_60;
output 	in_narrow_reg1;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Decoder1;
input 	Add2;
input 	Add21;
input 	Add22;
output 	nxt_out_eop;
input 	Equal2;
input 	src_valid;
input 	src_valid1;
output 	out_byte_cnt_reg_2;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	nxt_out_burstwrap_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \d0_int_bytes_remaining[2]~3_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[3]~4_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~0_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~1_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~2_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;


terminal_qsys_altera_merlin_address_alignment_5 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[79]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.src_payload2(sink0_data[78]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[60] (
	.clk(clk_clk),
	.d(sink0_data[60]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(!cp_ready),
	.datae(!\new_burst_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000004400000044;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!in_ready_hold),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'hA0A0F5F50000FF77;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!in_data_reg_60),
	.datad(!cp_ready),
	.datae(!\new_burst_reg~q ),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h0A0A0A4E5F1B5F5F;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(clk_clk),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(clk_clk),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(clk_clk),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(clk_clk),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(clk_clk),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(clk_clk),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[100] (
	.clk(clk_clk),
	.d(sink0_data[100]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_100),
	.prn(vcc));
defparam \in_data_reg[100] .is_wysiwyg = "true";
defparam \in_data_reg[100] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(clk_clk),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(clk_clk),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(clk_clk),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h0202020202020202;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0202020202020202;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h7777777777777777;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold),
	.datab(!nxt_out_eop),
	.datac(!src_valid),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h05CD05CD05CD05CD;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\Selector2~0_combout ),
	.datab(!in_data_reg_60),
	.datac(!nxt_out_eop),
	.datad(!src_valid),
	.datae(!stateST_COMP_TRANS),
	.dataf(!in_ready_hold),
	.datag(!\state.ST_IDLE~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "on";
defparam \Selector1~0 .lut_mask = 64'h0000F0F000F1F0FF;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!sink0_data[60]),
	.datab(!Equal2),
	.datac(!in_ready_hold),
	.datad(!nxt_in_ready),
	.datae(!nxt_in_ready1),
	.dataf(!src_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0000000001010001;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~3 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!sink0_data[60]),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~3 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~3 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~4 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!sink0_data[60]),
	.datad(!h2f_lw_ARLEN_1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_lw_ARLEN_0),
	.datag(!\int_bytes_remaining_reg[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~4 .extended_lut = "on";
defparam \d0_int_bytes_remaining[3]~4 .lut_mask = 64'h6363000F63630F00;
defparam \d0_int_bytes_remaining[3]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hA6AAA6AAA6AAA6AA;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~0 (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~0 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\int_bytes_remaining_reg[4]~q ),
	.datab(!\int_bytes_remaining_reg[3]~q ),
	.datac(!out_byte_cnt_reg_2),
	.datad(!\int_bytes_remaining_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0800080008000800;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~1 (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~1 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~2 (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~2 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\d0_int_bytes_remaining[4]~0_combout ),
	.datac(!\d0_int_bytes_remaining[5]~1_combout ),
	.datad(!\d0_int_bytes_remaining[6]~2_combout ),
	.datae(!\d0_int_bytes_remaining[2]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hAAAAEAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!sink0_data[60]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!mem_used_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0D8F0D8F0D8F0D8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_ready_hold),
	.datac(!src_valid),
	.datad(!\nxt_out_valid~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h0357035703570357;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h2020202020202020;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[73]),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\d0_int_nxt_addr[3]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[79]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[78]),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0044A0E40044A0E4;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[70]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[70]),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!sink0_data[60]),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!sink0_data[60]),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_lw_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!sink0_data[60]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!sink0_data[60]),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[72]),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\d0_int_nxt_addr[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!sink0_data[60]),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_address_alignment_5 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_2,
	src_payload2,
	in_size_reg_1,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_2;
input 	src_payload2;
input 	in_size_reg_1;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_2),
	.datad(!src_payload2),
	.datae(!in_size_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_adapter_5 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	Add5,
	Add51,
	Equal5,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_60,
	in_ready_hold,
	in_narrow_reg,
	cp_ready,
	nxt_in_ready,
	out_valid_reg,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	altera_reset_synchronizer_int_chain_out,
	nxt_out_eop,
	last_cycle,
	Decoder1,
	out_byte_cnt_reg_2,
	Add2,
	Add21,
	Add22,
	cp_ready1,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	Selector10,
	Selector101,
	Selector11,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add3,
	Selector12,
	Decoder11,
	src_payload,
	src_payload1,
	src_payload2,
	nxt_out_burstwrap_1,
	nxt_out_burstwrap_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	Add5;
input 	Add51;
input 	Equal5;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_60;
output 	in_ready_hold;
output 	in_narrow_reg;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	altera_reset_synchronizer_int_chain_out;
output 	nxt_out_eop;
input 	last_cycle;
input 	Decoder1;
output 	out_byte_cnt_reg_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	Selector10;
input 	Selector101;
input 	Selector11;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add3;
input 	Selector12;
input 	Decoder11;
input 	src_payload;
input 	src_payload1;
input 	src_payload2;
output 	nxt_out_burstwrap_1;
output 	nxt_out_burstwrap_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_adapter_13_1_5 \altera_merlin_burst_adapter_13_1.burst_adapter (
	.h2f_lw_ARADDR_0(h2f_lw_ARADDR_0),
	.h2f_lw_ARADDR_1(h2f_lw_ARADDR_1),
	.h2f_lw_ARADDR_2(h2f_lw_ARADDR_2),
	.h2f_lw_ARADDR_3(h2f_lw_ARADDR_3),
	.h2f_lw_ARBURST_0(h2f_lw_ARBURST_0),
	.h2f_lw_ARBURST_1(h2f_lw_ARBURST_1),
	.sink0_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,h2f_lw_ARID_11,h2f_lw_ARID_10,h2f_lw_ARID_9,h2f_lw_ARID_8,h2f_lw_ARID_7,h2f_lw_ARID_6,h2f_lw_ARID_5,h2f_lw_ARID_4,h2f_lw_ARID_3,h2f_lw_ARID_2,h2f_lw_ARID_1,h2f_lw_ARID_0,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload1,src_payload2,
src_payload,gnd,gnd,gnd,Selector101,Selector11,Selector12,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd}),
	.h2f_lw_ARLEN_0(h2f_lw_ARLEN_0),
	.h2f_lw_ARLEN_1(h2f_lw_ARLEN_1),
	.h2f_lw_ARLEN_2(h2f_lw_ARLEN_2),
	.h2f_lw_ARLEN_3(h2f_lw_ARLEN_3),
	.Add5(Add5),
	.Add51(Add51),
	.Equal5(Equal5),
	.saved_grant_1(saved_grant_1),
	.stateST_COMP_TRANS(stateST_COMP_TRANS),
	.mem_used_1(mem_used_1),
	.in_data_reg_60(in_data_reg_60),
	.in_ready_hold1(in_ready_hold),
	.in_narrow_reg1(in_narrow_reg),
	.cp_ready(cp_ready),
	.nxt_in_ready(nxt_in_ready),
	.out_valid_reg1(out_valid_reg),
	.stateST_UNCOMP_WR_SUBBURST(stateST_UNCOMP_WR_SUBBURST),
	.nxt_in_ready1(nxt_in_ready1),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.nxt_out_eop(nxt_out_eop),
	.last_cycle(last_cycle),
	.Decoder1(Decoder1),
	.out_byte_cnt_reg_2(out_byte_cnt_reg_2),
	.Add2(Add2),
	.Add21(Add21),
	.Add22(Add22),
	.cp_ready1(cp_ready1),
	.out_uncomp_byte_cnt_reg_5(out_uncomp_byte_cnt_reg_5),
	.out_uncomp_byte_cnt_reg_4(out_uncomp_byte_cnt_reg_4),
	.out_uncomp_byte_cnt_reg_3(out_uncomp_byte_cnt_reg_3),
	.out_uncomp_byte_cnt_reg_2(out_uncomp_byte_cnt_reg_2),
	.out_uncomp_byte_cnt_reg_6(out_uncomp_byte_cnt_reg_6),
	.in_data_reg_92(in_data_reg_92),
	.in_data_reg_93(in_data_reg_93),
	.in_data_reg_94(in_data_reg_94),
	.in_data_reg_95(in_data_reg_95),
	.in_data_reg_96(in_data_reg_96),
	.in_data_reg_97(in_data_reg_97),
	.in_data_reg_98(in_data_reg_98),
	.in_data_reg_99(in_data_reg_99),
	.in_data_reg_100(in_data_reg_100),
	.in_data_reg_101(in_data_reg_101),
	.in_data_reg_102(in_data_reg_102),
	.in_data_reg_103(in_data_reg_103),
	.Selector10(Selector10),
	.int_nxt_addr_reg_dly_3(int_nxt_addr_reg_dly_3),
	.int_nxt_addr_reg_dly_2(int_nxt_addr_reg_dly_2),
	.Add3(Add3),
	.Decoder11(Decoder11),
	.nxt_out_burstwrap_1(nxt_out_burstwrap_1),
	.nxt_out_burstwrap_0(nxt_out_burstwrap_0),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_merlin_burst_adapter_13_1_5 (
	h2f_lw_ARADDR_0,
	h2f_lw_ARADDR_1,
	h2f_lw_ARADDR_2,
	h2f_lw_ARADDR_3,
	h2f_lw_ARBURST_0,
	h2f_lw_ARBURST_1,
	sink0_data,
	h2f_lw_ARLEN_0,
	h2f_lw_ARLEN_1,
	h2f_lw_ARLEN_2,
	h2f_lw_ARLEN_3,
	Add5,
	Add51,
	Equal5,
	saved_grant_1,
	stateST_COMP_TRANS,
	mem_used_1,
	in_data_reg_60,
	in_ready_hold1,
	in_narrow_reg1,
	cp_ready,
	nxt_in_ready,
	out_valid_reg1,
	stateST_UNCOMP_WR_SUBBURST,
	nxt_in_ready1,
	altera_reset_synchronizer_int_chain_out,
	nxt_out_eop,
	last_cycle,
	Decoder1,
	out_byte_cnt_reg_2,
	Add2,
	Add21,
	Add22,
	cp_ready1,
	out_uncomp_byte_cnt_reg_5,
	out_uncomp_byte_cnt_reg_4,
	out_uncomp_byte_cnt_reg_3,
	out_uncomp_byte_cnt_reg_2,
	out_uncomp_byte_cnt_reg_6,
	in_data_reg_92,
	in_data_reg_93,
	in_data_reg_94,
	in_data_reg_95,
	in_data_reg_96,
	in_data_reg_97,
	in_data_reg_98,
	in_data_reg_99,
	in_data_reg_100,
	in_data_reg_101,
	in_data_reg_102,
	in_data_reg_103,
	Selector10,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	Add3,
	Decoder11,
	nxt_out_burstwrap_1,
	nxt_out_burstwrap_0,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_0;
input 	h2f_lw_ARADDR_1;
input 	h2f_lw_ARADDR_2;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARBURST_0;
input 	h2f_lw_ARBURST_1;
input 	[115:0] sink0_data;
input 	h2f_lw_ARLEN_0;
input 	h2f_lw_ARLEN_1;
input 	h2f_lw_ARLEN_2;
input 	h2f_lw_ARLEN_3;
input 	Add5;
input 	Add51;
input 	Equal5;
input 	saved_grant_1;
output 	stateST_COMP_TRANS;
input 	mem_used_1;
output 	in_data_reg_60;
output 	in_ready_hold1;
output 	in_narrow_reg1;
input 	cp_ready;
output 	nxt_in_ready;
output 	out_valid_reg1;
output 	stateST_UNCOMP_WR_SUBBURST;
output 	nxt_in_ready1;
input 	altera_reset_synchronizer_int_chain_out;
output 	nxt_out_eop;
input 	last_cycle;
input 	Decoder1;
output 	out_byte_cnt_reg_2;
input 	Add2;
input 	Add21;
input 	Add22;
input 	cp_ready1;
output 	out_uncomp_byte_cnt_reg_5;
output 	out_uncomp_byte_cnt_reg_4;
output 	out_uncomp_byte_cnt_reg_3;
output 	out_uncomp_byte_cnt_reg_2;
output 	out_uncomp_byte_cnt_reg_6;
output 	in_data_reg_92;
output 	in_data_reg_93;
output 	in_data_reg_94;
output 	in_data_reg_95;
output 	in_data_reg_96;
output 	in_data_reg_97;
output 	in_data_reg_98;
output 	in_data_reg_99;
output 	in_data_reg_100;
output 	in_data_reg_101;
output 	in_data_reg_102;
output 	in_data_reg_103;
input 	Selector10;
output 	int_nxt_addr_reg_dly_3;
output 	int_nxt_addr_reg_dly_2;
input 	Add3;
input 	Decoder11;
output 	nxt_out_burstwrap_1;
output 	nxt_out_burstwrap_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \align_address_to_size|LessThan0~0_combout ;
wire \align_address_to_size|LessThan0~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt~0_combout ;
wire \Add4~0_combout ;
wire \nxt_uncomp_subburst_byte_cnt[5]~1_combout ;
wire \nxt_uncomp_subburst_byte_cnt[6]~2_combout ;
wire \nxt_uncomp_subburst_byte_cnt[3]~3_combout ;
wire \nxt_uncomp_subburst_byte_cnt[4]~4_combout ;
wire \nxt_uncomp_subburst_byte_cnt[2]~5_combout ;
wire \WideNor1~combout ;
wire \Selector2~1_combout ;
wire \load_next_out_cmd~combout ;
wire \state.ST_UNCOMP_TRANS~q ;
wire \Selector2~0_combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \NON_PIPELINED_INPUTS.load_next_cmd~0_combout ;
wire \int_bytes_remaining_reg[2]~q ;
wire \d0_int_bytes_remaining[2]~0_combout ;
wire \int_bytes_remaining_reg[4]~q ;
wire \d0_int_bytes_remaining[3]~4_combout ;
wire \int_bytes_remaining_reg[3]~q ;
wire \Add1~0_combout ;
wire \d0_int_bytes_remaining[4]~1_combout ;
wire \int_bytes_remaining_reg[5]~q ;
wire \Add1~1_combout ;
wire \d0_int_bytes_remaining[5]~2_combout ;
wire \int_bytes_remaining_reg[6]~q ;
wire \d0_int_bytes_remaining[6]~3_combout ;
wire \new_burst_reg~0_combout ;
wire \new_burst_reg~q ;
wire \in_bytecount_reg_zero~0_combout ;
wire \in_bytecount_reg_zero~q ;
wire \nxt_out_valid~0_combout ;
wire \nxt_out_valid~1_combout ;
wire \Selector3~0_combout ;
wire \in_burstwrap_reg[3]~q ;
wire \nxt_addr[3]~combout ;
wire \int_nxt_addr_reg[3]~q ;
wire \in_size_reg[0]~q ;
wire \in_size_reg[2]~q ;
wire \in_size_reg[1]~q ;
wire \ShiftLeft0~0_combout ;
wire \ShiftLeft0~1_combout ;
wire \int_byte_cnt_narrow_reg[3]~q ;
wire \ShiftLeft0~2_combout ;
wire \int_byte_cnt_narrow_reg[2]~q ;
wire \in_burstwrap_reg[1]~q ;
wire \nxt_addr[1]~combout ;
wire \int_nxt_addr_reg[1]~q ;
wire \ShiftLeft0~3_combout ;
wire \int_byte_cnt_narrow_reg[1]~q ;
wire \int_byte_cnt_narrow_reg[0]~q ;
wire \Add0~13_sumout ;
wire \in_burstwrap_reg[0]~q ;
wire \nxt_addr[0]~combout ;
wire \int_nxt_addr_reg[0]~q ;
wire \d0_int_nxt_addr[0]~2_combout ;
wire \d0_int_nxt_addr[0]~3_combout ;
wire \int_nxt_addr_reg_dly[0]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \d0_int_nxt_addr[1]~4_combout ;
wire \int_nxt_addr_reg_dly[1]~q ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \d0_int_nxt_addr[3]~0_combout ;
wire \in_burstwrap_reg[2]~q ;
wire \nxt_addr[2]~combout ;
wire \int_nxt_addr_reg[2]~q ;
wire \Add0~5_sumout ;
wire \d0_int_nxt_addr[2]~1_combout ;
wire \nxt_out_burstwrap[0]~1_combout ;


terminal_qsys_altera_merlin_address_alignment_6 align_address_to_size(
	.new_burst_reg(\new_burst_reg~q ),
	.src_payload(sink0_data[77]),
	.in_size_reg_0(\in_size_reg[0]~q ),
	.src_payload1(sink0_data[79]),
	.in_size_reg_2(\in_size_reg[2]~q ),
	.src_payload2(sink0_data[78]),
	.in_size_reg_1(\in_size_reg[1]~q ),
	.LessThan0(\align_address_to_size|LessThan0~0_combout ),
	.LessThan01(\align_address_to_size|LessThan0~1_combout ));

dffeas \state.ST_COMP_TRANS (
	.clk(clk_clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_COMP_TRANS),
	.prn(vcc));
defparam \state.ST_COMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_COMP_TRANS .power_up = "low";

dffeas \in_data_reg[60] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_60),
	.prn(vcc));
defparam \in_data_reg[60] .is_wysiwyg = "true";
defparam \in_data_reg[60] .power_up = "low";

dffeas in_ready_hold(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_hold1),
	.prn(vcc));
defparam in_ready_hold.is_wysiwyg = "true";
defparam in_ready_hold.power_up = "low";

dffeas in_narrow_reg(
	.clk(clk_clk),
	.d(Decoder1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_narrow_reg1),
	.prn(vcc));
defparam in_narrow_reg.is_wysiwyg = "true";
defparam in_narrow_reg.power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(!cp_ready),
	.datae(!\new_burst_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~0 .extended_lut = "off";
defparam \nxt_in_ready~0 .lut_mask = 64'h0000004400000044;
defparam \nxt_in_ready~0 .shared_arith = "off";

dffeas out_valid_reg(
	.clk(clk_clk),
	.d(\nxt_out_valid~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_valid_reg1),
	.prn(vcc));
defparam out_valid_reg.is_wysiwyg = "true";
defparam out_valid_reg.power_up = "low";

dffeas \state.ST_UNCOMP_WR_SUBBURST (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(stateST_UNCOMP_WR_SUBBURST),
	.prn(vcc));
defparam \state.ST_UNCOMP_WR_SUBBURST .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_WR_SUBBURST .power_up = "low";

cyclonev_lcell_comb \nxt_in_ready~1 (
	.dataa(!in_ready_hold1),
	.datab(!stateST_COMP_TRANS),
	.datac(!mem_used_1),
	.datad(!cp_ready),
	.datae(!out_valid_reg1),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_in_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_in_ready~1 .extended_lut = "off";
defparam \nxt_in_ready~1 .lut_mask = 64'h0000FF3F8888BBBB;
defparam \nxt_in_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_eop~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!mem_used_1),
	.datac(!in_data_reg_60),
	.datad(!cp_ready),
	.datae(!\new_burst_reg~q ),
	.dataf(!\in_bytecount_reg_zero~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_eop),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_eop~0 .extended_lut = "off";
defparam \nxt_out_eop~0 .lut_mask = 64'h0A0A0A4E5F1B5F5F;
defparam \nxt_out_eop~0 .shared_arith = "off";

dffeas \out_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[5] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_5),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[5] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[5] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[4] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_4),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[4] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[4] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[3] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_3),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[3] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[3] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[2] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_2),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[2] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[2] .power_up = "low";

dffeas \out_uncomp_byte_cnt_reg[6] (
	.clk(clk_clk),
	.d(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(out_uncomp_byte_cnt_reg_6),
	.prn(vcc));
defparam \out_uncomp_byte_cnt_reg[6] .is_wysiwyg = "true";
defparam \out_uncomp_byte_cnt_reg[6] .power_up = "low";

dffeas \in_data_reg[92] (
	.clk(clk_clk),
	.d(sink0_data[92]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_92),
	.prn(vcc));
defparam \in_data_reg[92] .is_wysiwyg = "true";
defparam \in_data_reg[92] .power_up = "low";

dffeas \in_data_reg[93] (
	.clk(clk_clk),
	.d(sink0_data[93]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_93),
	.prn(vcc));
defparam \in_data_reg[93] .is_wysiwyg = "true";
defparam \in_data_reg[93] .power_up = "low";

dffeas \in_data_reg[94] (
	.clk(clk_clk),
	.d(sink0_data[94]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_94),
	.prn(vcc));
defparam \in_data_reg[94] .is_wysiwyg = "true";
defparam \in_data_reg[94] .power_up = "low";

dffeas \in_data_reg[95] (
	.clk(clk_clk),
	.d(sink0_data[95]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_95),
	.prn(vcc));
defparam \in_data_reg[95] .is_wysiwyg = "true";
defparam \in_data_reg[95] .power_up = "low";

dffeas \in_data_reg[96] (
	.clk(clk_clk),
	.d(sink0_data[96]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_96),
	.prn(vcc));
defparam \in_data_reg[96] .is_wysiwyg = "true";
defparam \in_data_reg[96] .power_up = "low";

dffeas \in_data_reg[97] (
	.clk(clk_clk),
	.d(sink0_data[97]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_97),
	.prn(vcc));
defparam \in_data_reg[97] .is_wysiwyg = "true";
defparam \in_data_reg[97] .power_up = "low";

dffeas \in_data_reg[98] (
	.clk(clk_clk),
	.d(sink0_data[98]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_98),
	.prn(vcc));
defparam \in_data_reg[98] .is_wysiwyg = "true";
defparam \in_data_reg[98] .power_up = "low";

dffeas \in_data_reg[99] (
	.clk(clk_clk),
	.d(sink0_data[99]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_99),
	.prn(vcc));
defparam \in_data_reg[99] .is_wysiwyg = "true";
defparam \in_data_reg[99] .power_up = "low";

dffeas \in_data_reg[100] (
	.clk(clk_clk),
	.d(sink0_data[100]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_100),
	.prn(vcc));
defparam \in_data_reg[100] .is_wysiwyg = "true";
defparam \in_data_reg[100] .power_up = "low";

dffeas \in_data_reg[101] (
	.clk(clk_clk),
	.d(sink0_data[101]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_101),
	.prn(vcc));
defparam \in_data_reg[101] .is_wysiwyg = "true";
defparam \in_data_reg[101] .power_up = "low";

dffeas \in_data_reg[102] (
	.clk(clk_clk),
	.d(sink0_data[102]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_102),
	.prn(vcc));
defparam \in_data_reg[102] .is_wysiwyg = "true";
defparam \in_data_reg[102] .power_up = "low";

dffeas \in_data_reg[103] (
	.clk(clk_clk),
	.d(sink0_data[103]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(in_data_reg_103),
	.prn(vcc));
defparam \in_data_reg[103] .is_wysiwyg = "true";
defparam \in_data_reg[103] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[3] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_3),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[3] .power_up = "low";

dffeas \int_nxt_addr_reg_dly[2] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(int_nxt_addr_reg_dly_2),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[2] .power_up = "low";

cyclonev_lcell_comb \nxt_out_burstwrap[1]~0 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!Selector10),
	.datad(!Add3),
	.datae(!Add5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_burstwrap_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[1]~0 .extended_lut = "off";
defparam \nxt_out_burstwrap[1]~0 .lut_mask = 64'h8A8802008A880200;
defparam \nxt_out_burstwrap[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_burstwrap[0]~2 (
	.dataa(!h2f_lw_ARBURST_0),
	.datab(!h2f_lw_ARBURST_1),
	.datac(!Decoder11),
	.datad(!Add51),
	.datae(!\nxt_out_burstwrap[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nxt_out_burstwrap_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[0]~2 .extended_lut = "off";
defparam \nxt_out_burstwrap[0]~2 .lut_mask = 64'h77FF75FD77FF75FD;
defparam \nxt_out_burstwrap[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt~0 (
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt~0 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt~0 .lut_mask = 64'h0202020202020202;
defparam \nxt_uncomp_subburst_byte_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!out_uncomp_byte_cnt_reg_4),
	.datab(!out_uncomp_byte_cnt_reg_3),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h0800080008000800;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[5]~1 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .lut_mask = 64'h0F4EA5E40F4EA5E4;
defparam \nxt_uncomp_subburst_byte_cnt[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[6]~2 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_5),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!\Add4~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .lut_mask = 64'h0044A0E4FFEE5F4E;
defparam \nxt_uncomp_subburst_byte_cnt[6]~2 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[3]~3 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_3),
	.datad(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datae(!out_uncomp_byte_cnt_reg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .lut_mask = 64'h0FE40F4E0FE40F4E;
defparam \nxt_uncomp_subburst_byte_cnt[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[4]~4 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!out_uncomp_byte_cnt_reg_4),
	.datad(!out_uncomp_byte_cnt_reg_3),
	.datae(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.dataf(!out_uncomp_byte_cnt_reg_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .lut_mask = 64'h0F0FE44E0F0F4E4E;
defparam \nxt_uncomp_subburst_byte_cnt[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \nxt_uncomp_subburst_byte_cnt[2]~5 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!\nxt_uncomp_subburst_byte_cnt~0_combout ),
	.datad(!out_uncomp_byte_cnt_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .extended_lut = "off";
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .lut_mask = 64'h0EF40EF40EF40EF4;
defparam \nxt_uncomp_subburst_byte_cnt[2]~5 .shared_arith = "off";

cyclonev_lcell_comb WideNor1(
	.dataa(!\nxt_uncomp_subburst_byte_cnt[5]~1_combout ),
	.datab(!\nxt_uncomp_subburst_byte_cnt[6]~2_combout ),
	.datac(!\nxt_uncomp_subburst_byte_cnt[3]~3_combout ),
	.datad(!\nxt_uncomp_subburst_byte_cnt[4]~4_combout ),
	.datae(!\nxt_uncomp_subburst_byte_cnt[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h8000000080000000;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h0808080808080808;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb load_next_out_cmd(
	.dataa(!mem_used_1),
	.datab(!cp_ready),
	.datac(!out_valid_reg1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_next_out_cmd~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam load_next_out_cmd.extended_lut = "off";
defparam load_next_out_cmd.lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam load_next_out_cmd.shared_arith = "off";

dffeas \state.ST_UNCOMP_TRANS (
	.clk(clk_clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_UNCOMP_TRANS~q ),
	.prn(vcc));
defparam \state.ST_UNCOMP_TRANS .is_wysiwyg = "true";
defparam \state.ST_UNCOMP_TRANS .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\state.ST_UNCOMP_TRANS~q ),
	.datab(!stateST_UNCOMP_WR_SUBBURST),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h8888888888888888;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!in_ready_hold1),
	.datab(!Equal5),
	.datac(!nxt_out_eop),
	.datad(!last_cycle),
	.datae(!\state.ST_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h0011F0F10011F0F1;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_data_reg_60),
	.datac(!\Selector2~0_combout ),
	.datad(!\state.ST_IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h008A008A008A008A;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!in_ready_hold1),
	.datab(!Equal5),
	.datac(!stateST_COMP_TRANS),
	.datad(!nxt_out_eop),
	.datae(!last_cycle),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h0F001F110F000F00;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \NON_PIPELINED_INPUTS.load_next_cmd~0 (
	.dataa(!in_ready_hold1),
	.datab(!Equal5),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(!last_cycle),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .extended_lut = "off";
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .lut_mask = 64'h0000110100001101;
defparam \NON_PIPELINED_INPUTS.load_next_cmd~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[2] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[2]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[2]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[2] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[2]~0 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!out_byte_cnt_reg_2),
	.datae(!\int_bytes_remaining_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[2]~0 .extended_lut = "off";
defparam \d0_int_bytes_remaining[2]~0 .lut_mask = 64'h02F2F20202F2F202;
defparam \d0_int_bytes_remaining[2]~0 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[4] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[4]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[4] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[4] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[3]~4 (
	.dataa(!\int_bytes_remaining_reg[2]~q ),
	.datab(!out_byte_cnt_reg_2),
	.datac(!saved_grant_1),
	.datad(!h2f_lw_ARLEN_1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_lw_ARLEN_0),
	.datag(!\int_bytes_remaining_reg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[3]~4 .extended_lut = "on";
defparam \d0_int_bytes_remaining[3]~4 .lut_mask = 64'h2D2D000F2D2D0F00;
defparam \d0_int_bytes_remaining[3]~4 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[3] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[3]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[3] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[3] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hB4F0B4F0B4F0B4F0;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[4]~1 (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!Add2),
	.datad(!\Add1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[4]~1 .extended_lut = "off";
defparam \d0_int_bytes_remaining[4]~1 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \d0_int_bytes_remaining[4]~1 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[5] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[5]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[5] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!out_byte_cnt_reg_2),
	.datab(!\int_bytes_remaining_reg[2]~q ),
	.datac(!\int_bytes_remaining_reg[4]~q ),
	.datad(!\int_bytes_remaining_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h4000400040004000;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_bytes_remaining[5]~2 (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!Add21),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[5]~2 .extended_lut = "off";
defparam \d0_int_bytes_remaining[5]~2 .lut_mask = 64'h01CDCD0101CDCD01;
defparam \d0_int_bytes_remaining[5]~2 .shared_arith = "off";

dffeas \int_bytes_remaining_reg[6] (
	.clk(clk_clk),
	.d(\d0_int_bytes_remaining[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_bytes_remaining_reg[6]~q ),
	.prn(vcc));
defparam \int_bytes_remaining_reg[6] .is_wysiwyg = "true";
defparam \int_bytes_remaining_reg[6] .power_up = "low";

cyclonev_lcell_comb \d0_int_bytes_remaining[6]~3 (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!Add22),
	.datad(!\int_bytes_remaining_reg[5]~q ),
	.datae(!\Add1~1_combout ),
	.dataf(!\int_bytes_remaining_reg[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_bytes_remaining[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_bytes_remaining[6]~3 .extended_lut = "off";
defparam \d0_int_bytes_remaining[6]~3 .lut_mask = 64'h0101CD01CDCD01CD;
defparam \d0_int_bytes_remaining[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \new_burst_reg~0 (
	.dataa(!\Selector1~1_combout ),
	.datab(!\d0_int_bytes_remaining[2]~0_combout ),
	.datac(!\d0_int_bytes_remaining[4]~1_combout ),
	.datad(!\d0_int_bytes_remaining[5]~2_combout ),
	.datae(!\d0_int_bytes_remaining[6]~3_combout ),
	.dataf(!\d0_int_bytes_remaining[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_burst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_burst_reg~0 .extended_lut = "off";
defparam \new_burst_reg~0 .lut_mask = 64'hBAAAAAAAAAAAAAAA;
defparam \new_burst_reg~0 .shared_arith = "off";

dffeas new_burst_reg(
	.clk(clk_clk),
	.d(\new_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\new_burst_reg~q ),
	.prn(vcc));
defparam new_burst_reg.is_wysiwyg = "true";
defparam new_burst_reg.power_up = "low";

cyclonev_lcell_comb \in_bytecount_reg_zero~0 (
	.dataa(!saved_grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\in_bytecount_reg_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \in_bytecount_reg_zero~0 .extended_lut = "off";
defparam \in_bytecount_reg_zero~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \in_bytecount_reg_zero~0 .shared_arith = "off";

dffeas in_bytecount_reg_zero(
	.clk(clk_clk),
	.d(\in_bytecount_reg_zero~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_bytecount_reg_zero~q ),
	.prn(vcc));
defparam in_bytecount_reg_zero.is_wysiwyg = "true";
defparam in_bytecount_reg_zero.power_up = "low";

cyclonev_lcell_comb \nxt_out_valid~0 (
	.dataa(!mem_used_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_bytecount_reg_zero~q ),
	.datad(!cp_ready1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~0 .extended_lut = "off";
defparam \nxt_out_valid~0 .lut_mask = 64'hF0D8F0D8F0D8F0D8;
defparam \nxt_out_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_valid~1 (
	.dataa(!in_ready_hold1),
	.datab(!Equal5),
	.datac(!stateST_COMP_TRANS),
	.datad(!last_cycle),
	.datae(!\nxt_out_valid~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_valid~1 .extended_lut = "off";
defparam \nxt_out_valid~1 .lut_mask = 64'h00110F1F00110F1F;
defparam \nxt_out_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!nxt_out_eop),
	.datab(!\Selector2~0_combout ),
	.datac(!\WideNor1~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h8080808080808080;
defparam \Selector3~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[3] (
	.clk(clk_clk),
	.d(sink0_data[73]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[3]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[3] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[3] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[3] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[73]),
	.datad(!\in_burstwrap_reg[3]~q ),
	.datae(!\d0_int_nxt_addr[3]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[3] .extended_lut = "off";
defparam \nxt_addr[3] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[3] .shared_arith = "off";

dffeas \int_nxt_addr_reg[3] (
	.clk(clk_clk),
	.d(\nxt_addr[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[3]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[3] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[3] .power_up = "low";

dffeas \in_size_reg[0] (
	.clk(clk_clk),
	.d(sink0_data[77]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[0]~q ),
	.prn(vcc));
defparam \in_size_reg[0] .is_wysiwyg = "true";
defparam \in_size_reg[0] .power_up = "low";

dffeas \in_size_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[79]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[2]~q ),
	.prn(vcc));
defparam \in_size_reg[2] .is_wysiwyg = "true";
defparam \in_size_reg[2] .power_up = "low";

dffeas \in_size_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[78]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_size_reg[1]~q ),
	.prn(vcc));
defparam \in_size_reg[1] .is_wysiwyg = "true";
defparam \in_size_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~0 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[79]),
	.datac(!\in_size_reg[2]~q ),
	.datad(!sink0_data[78]),
	.datae(!\in_size_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~0 .extended_lut = "off";
defparam \ShiftLeft0~0 .lut_mask = 64'h0044A0E40044A0E4;
defparam \ShiftLeft0~0 .shared_arith = "off";

cyclonev_lcell_comb \ShiftLeft0~1 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~1 .extended_lut = "off";
defparam \ShiftLeft0~1 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~1 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[3] (
	.clk(clk_clk),
	.d(\ShiftLeft0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[3]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[3] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[3] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~2 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\ShiftLeft0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~2 .extended_lut = "off";
defparam \ShiftLeft0~2 .lut_mask = 64'h00E400E400E400E4;
defparam \ShiftLeft0~2 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[2] (
	.clk(clk_clk),
	.d(\ShiftLeft0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[2]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[2] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[2] .power_up = "low";

dffeas \in_burstwrap_reg[1] (
	.clk(clk_clk),
	.d(sink0_data[71]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[1]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[1] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[1] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[1] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!\in_burstwrap_reg[1]~q ),
	.datad(!\d0_int_nxt_addr[1]~4_combout ),
	.datae(!nxt_out_burstwrap_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[1] .extended_lut = "off";
defparam \nxt_addr[1] .lut_mask = 64'h00E200F300E200F3;
defparam \nxt_addr[1] .shared_arith = "off";

dffeas \int_nxt_addr_reg[1] (
	.clk(clk_clk),
	.d(\nxt_addr[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[1] .power_up = "low";

cyclonev_lcell_comb \ShiftLeft0~3 (
	.dataa(!\new_burst_reg~q ),
	.datab(!sink0_data[77]),
	.datac(!\in_size_reg[0]~q ),
	.datad(!\align_address_to_size|LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ShiftLeft0~3 .extended_lut = "off";
defparam \ShiftLeft0~3 .lut_mask = 64'h001B001B001B001B;
defparam \ShiftLeft0~3 .shared_arith = "off";

dffeas \int_byte_cnt_narrow_reg[1] (
	.clk(clk_clk),
	.d(\ShiftLeft0~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[1]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[1] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[1] .power_up = "low";

dffeas \int_byte_cnt_narrow_reg[0] (
	.clk(clk_clk),
	.d(\align_address_to_size|LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_byte_cnt_narrow_reg[0]~q ),
	.prn(vcc));
defparam \int_byte_cnt_narrow_reg[0] .is_wysiwyg = "true";
defparam \int_byte_cnt_narrow_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[0]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \in_burstwrap_reg[0] (
	.clk(clk_clk),
	.d(nxt_out_burstwrap_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[0]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[0] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[0] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[0] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!nxt_out_burstwrap_0),
	.datad(!\in_burstwrap_reg[0]~q ),
	.datae(!\d0_int_nxt_addr[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[0] .extended_lut = "off";
defparam \nxt_addr[0] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[0] .shared_arith = "off";

dffeas \int_nxt_addr_reg[0] (
	.clk(clk_clk),
	.d(\nxt_addr[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[0] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~2 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\int_nxt_addr_reg[0]~q ),
	.datac(!\in_burstwrap_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~2 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~2 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \d0_int_nxt_addr[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[0]~3 (
	.dataa(!h2f_lw_ARADDR_0),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\align_address_to_size|LessThan0~1_combout ),
	.datae(!\d0_int_nxt_addr[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[0]~3 .extended_lut = "off";
defparam \d0_int_nxt_addr[0]~3 .lut_mask = 64'hF0F10001F0F10001;
defparam \d0_int_nxt_addr[0]~3 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[0] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[0]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[0] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\int_nxt_addr_reg_dly[1]~q ),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[1]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[1]~4 (
	.dataa(!\int_nxt_addr_reg[1]~q ),
	.datab(!\Add0~9_sumout ),
	.datac(!saved_grant_1),
	.datad(!Decoder1),
	.datae(!\new_burst_reg~q ),
	.dataf(!h2f_lw_ARADDR_1),
	.datag(!\in_burstwrap_reg[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[1]~4 .extended_lut = "on";
defparam \d0_int_nxt_addr[1]~4 .lut_mask = 64'h575700005757000F;
defparam \d0_int_nxt_addr[1]~4 .shared_arith = "off";

dffeas \int_nxt_addr_reg_dly[1] (
	.clk(clk_clk),
	.d(\d0_int_nxt_addr[1]~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg_dly[1]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg_dly[1] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg_dly[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_2),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[2]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!int_nxt_addr_reg_dly_3),
	.datae(gnd),
	.dataf(!\int_byte_cnt_narrow_reg[3]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \d0_int_nxt_addr[3]~0 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[3]~q ),
	.datae(!\in_burstwrap_reg[3]~q ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[3]~0 .extended_lut = "off";
defparam \d0_int_nxt_addr[3]~0 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[3]~0 .shared_arith = "off";

dffeas \in_burstwrap_reg[2] (
	.clk(clk_clk),
	.d(sink0_data[72]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\NON_PIPELINED_INPUTS.load_next_cmd~0_combout ),
	.q(\in_burstwrap_reg[2]~q ),
	.prn(vcc));
defparam \in_burstwrap_reg[2] .is_wysiwyg = "true";
defparam \in_burstwrap_reg[2] .power_up = "low";

cyclonev_lcell_comb \nxt_addr[2] (
	.dataa(!saved_grant_1),
	.datab(!\new_burst_reg~q ),
	.datac(!sink0_data[72]),
	.datad(!\in_burstwrap_reg[2]~q ),
	.datae(!\d0_int_nxt_addr[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_addr[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_addr[2] .extended_lut = "off";
defparam \nxt_addr[2] .lut_mask = 64'h0000FE320000FE32;
defparam \nxt_addr[2] .shared_arith = "off";

dffeas \int_nxt_addr_reg[2] (
	.clk(clk_clk),
	.d(\nxt_addr[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_next_out_cmd~combout ),
	.q(\int_nxt_addr_reg[2]~q ),
	.prn(vcc));
defparam \int_nxt_addr_reg[2] .is_wysiwyg = "true";
defparam \int_nxt_addr_reg[2] .power_up = "low";

cyclonev_lcell_comb \d0_int_nxt_addr[2]~1 (
	.dataa(!h2f_lw_ARADDR_2),
	.datab(!saved_grant_1),
	.datac(!\new_burst_reg~q ),
	.datad(!\int_nxt_addr_reg[2]~q ),
	.datae(!\in_burstwrap_reg[2]~q ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d0_int_nxt_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d0_int_nxt_addr[2]~1 .extended_lut = "off";
defparam \d0_int_nxt_addr[2]~1 .lut_mask = 64'h01F101F101F1F1F1;
defparam \d0_int_nxt_addr[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \nxt_out_burstwrap[0]~1 (
	.dataa(!h2f_lw_ARLEN_0),
	.datab(!h2f_lw_ARLEN_1),
	.datac(!h2f_lw_ARLEN_2),
	.datad(!h2f_lw_ARLEN_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nxt_out_burstwrap[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nxt_out_burstwrap[0]~1 .extended_lut = "off";
defparam \nxt_out_burstwrap[0]~1 .lut_mask = 64'h8000800080008000;
defparam \nxt_out_burstwrap[0]~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_address_alignment_6 (
	new_burst_reg,
	src_payload,
	in_size_reg_0,
	src_payload1,
	in_size_reg_2,
	src_payload2,
	in_size_reg_1,
	LessThan0,
	LessThan01)/* synthesis synthesis_greybox=0 */;
input 	new_burst_reg;
input 	src_payload;
input 	in_size_reg_0;
input 	src_payload1;
input 	in_size_reg_2;
input 	src_payload2;
input 	in_size_reg_1;
output 	LessThan0;
output 	LessThan01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!new_burst_reg),
	.datab(!src_payload1),
	.datac(!in_size_reg_2),
	.datad(!src_payload2),
	.datae(!in_size_reg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hE4A04400E4A04400;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!new_burst_reg),
	.datab(!src_payload),
	.datac(!in_size_reg_0),
	.datad(!LessThan0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan01),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h00E400E400E400E4;
defparam \LessThan0~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_slave_agent (
	stateST_COMP_TRANS,
	out_valid_reg,
	in_ready_hold,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_59,
	local_write1,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	mem_57_0,
	comb,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	cp_ready,
	last_packet_beat2,
	read,
	rp_valid1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	in_ready_hold;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
output 	local_write1;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	mem_57_0;
output 	comb;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
output 	cp_ready;
output 	last_packet_beat2;
input 	read;
output 	rp_valid1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~0_combout ;
wire \cp_ready~1_combout ;


terminal_qsys_altera_merlin_burst_uncompressor uncompressor(
	.mem_57_0(mem_57_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_59),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(local_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!local_write1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~0_combout ),
	.datad(!\cp_ready~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!local_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_uncompressor (
	mem_57_0,
	comb,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_57_0;
input 	comb;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_slave_agent_1 (
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_59,
	local_write1,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	mem_57_0,
	comb,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	cp_ready,
	last_packet_beat2,
	read,
	rp_valid1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
output 	local_write1;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	mem_57_0;
output 	comb;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
output 	cp_ready;
output 	last_packet_beat2;
input 	read;
output 	rp_valid1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cp_ready~0_combout ;
wire \cp_ready~1_combout ;


terminal_qsys_altera_merlin_burst_uncompressor_1 uncompressor(
	.mem_57_0(mem_57_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_59),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(local_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!local_write1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~2 (
	.dataa(!mem_used_1),
	.datab(!in_narrow_reg),
	.datac(!\cp_ready~0_combout ),
	.datad(!\cp_ready~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~2 .extended_lut = "off";
defparam \cp_ready~2 .lut_mask = 64'h08AA08AA08AA08AA;
defparam \cp_ready~2 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_byteen_reg_3),
	.datab(!in_byteen_reg_2),
	.datac(!in_byteen_reg_1),
	.datad(!in_byteen_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h8000800080008000;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!local_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cp_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_uncompressor_1 (
	mem_57_0,
	comb,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_57_0;
input 	comb;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_slave_agent_2 (
	in_ready_hold,
	stateST_COMP_TRANS,
	out_valid_reg,
	mem_used_1,
	in_narrow_reg,
	in_byteen_reg_3,
	in_byteen_reg_2,
	in_byteen_reg_1,
	in_byteen_reg_0,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	in_data_reg_59,
	local_write1,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	mem_57_0,
	comb,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	m0_write1,
	cp_ready,
	cp_ready1,
	last_packet_beat2,
	read,
	rp_valid1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	stateST_COMP_TRANS;
input 	out_valid_reg;
input 	mem_used_1;
input 	in_narrow_reg;
input 	in_byteen_reg_3;
input 	in_byteen_reg_2;
input 	in_byteen_reg_1;
input 	in_byteen_reg_0;
output 	WideOr0;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	in_data_reg_59;
output 	local_write1;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	mem_57_0;
output 	comb;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	m0_write1;
output 	cp_ready;
output 	cp_ready1;
output 	last_packet_beat2;
input 	read;
output 	rp_valid1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_uncompressor_2 uncompressor(
	.mem_57_0(mem_57_0),
	.comb(comb),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_narrow_reg),
	.datac(!in_byteen_reg_3),
	.datad(!in_byteen_reg_2),
	.datae(!in_byteen_reg_1),
	.dataf(!in_byteen_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h1FFFFFFFFFFFFFFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb local_write(
	.dataa(!in_data_reg_59),
	.datab(!out_valid_reg),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(local_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam local_write.extended_lut = "off";
defparam local_write.lut_mask = 64'h1111111111111111;
defparam local_write.shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h007F007F007F007F;
defparam \comb~0 .shared_arith = "off";

cyclonev_lcell_comb m0_write(
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!local_write1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam m0_write.extended_lut = "off";
defparam m0_write.lut_mask = 64'h0202020202020202;
defparam m0_write.shared_arith = "off";

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_narrow_reg),
	.datab(!in_byteen_reg_3),
	.datac(!in_byteen_reg_2),
	.datad(!in_byteen_reg_1),
	.datae(!in_byteen_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'h8000000080000000;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!local_write1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h0440044004400440;
defparam \cp_ready~1 .shared_arith = "off";

cyclonev_lcell_comb rp_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rp_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam rp_valid.extended_lut = "off";
defparam rp_valid.lut_mask = 64'h8880888088808880;
defparam rp_valid.shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_uncompressor_2 (
	mem_57_0,
	comb,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	mem_57_0;
input 	comb;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!last_packet_beat),
	.datad(!last_packet_beat1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3222322232223222;
defparam \last_packet_beat~2 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(read),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_slave_agent_3 (
	in_ready_hold,
	stateST_COMP_TRANS,
	in_data_reg_60,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	empty,
	mem_57_0,
	mem_used_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	read,
	cp_ready1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	stateST_COMP_TRANS;
input 	in_data_reg_60;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
input 	empty;
input 	mem_57_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
input 	read;
output 	cp_ready1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_uncompressor_3 uncompressor(
	.empty(empty),
	.mem_57_0(mem_57_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_data_reg_60),
	.datac(!in_narrow_reg),
	.datad(!in_ready_hold),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC8C8C8C8C8FFC8C8;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_data_reg_60),
	.datab(!in_narrow_reg),
	.datac(!in_ready_hold),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h88888F8888888F88;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_uncompressor_3 (
	empty,
	mem_57_0,
	mem_used_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	empty;
input 	mem_57_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_57_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h1111111111111111;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_slave_agent_4 (
	in_ready_hold,
	stateST_COMP_TRANS,
	in_data_reg_60,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	empty,
	mem_57_0,
	mem_used_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	read,
	cp_ready1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	stateST_COMP_TRANS;
input 	in_data_reg_60;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
input 	empty;
input 	mem_57_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
input 	read;
output 	cp_ready1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_uncompressor_4 uncompressor(
	.empty(empty),
	.mem_57_0(mem_57_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!stateST_COMP_TRANS),
	.datab(!in_data_reg_60),
	.datac(!in_narrow_reg),
	.datad(!in_ready_hold),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hC8C8C8C8C8FFC8C8;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_data_reg_60),
	.datab(!in_narrow_reg),
	.datac(!in_ready_hold),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'h88888F8888888F88;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_uncompressor_4 (
	empty,
	mem_57_0,
	mem_used_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	empty;
input 	mem_57_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_57_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h1111111111111111;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_slave_agent_5 (
	stateST_COMP_TRANS,
	in_data_reg_60,
	in_ready_hold,
	in_narrow_reg,
	wait_latency_counter_1,
	wait_latency_counter_0,
	cp_ready,
	empty,
	mem_57_0,
	mem_used_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	altera_reset_synchronizer_int_chain_out,
	last_packet_beat2,
	read,
	cp_ready1,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	stateST_COMP_TRANS;
input 	in_data_reg_60;
input 	in_ready_hold;
input 	in_narrow_reg;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	cp_ready;
input 	empty;
input 	mem_57_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	altera_reset_synchronizer_int_chain_out;
output 	last_packet_beat2;
input 	read;
output 	cp_ready1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_merlin_burst_uncompressor_5 uncompressor(
	.empty(empty),
	.mem_57_0(mem_57_0),
	.mem_used_0(mem_used_0),
	.last_packet_beat(last_packet_beat),
	.mem_69_0(mem_69_0),
	.mem_68_0(mem_68_0),
	.mem_67_0(mem_67_0),
	.mem_66_0(mem_66_0),
	.mem_65_0(mem_65_0),
	.last_packet_beat1(last_packet_beat1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.last_packet_beat2(last_packet_beat2),
	.read(read),
	.clk(clk_clk));

cyclonev_lcell_comb \cp_ready~0 (
	.dataa(!in_ready_hold),
	.datab(!stateST_COMP_TRANS),
	.datac(!in_data_reg_60),
	.datad(!in_narrow_reg),
	.datae(!wait_latency_counter_1),
	.dataf(!wait_latency_counter_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~0 .extended_lut = "off";
defparam \cp_ready~0 .lut_mask = 64'hF0C0F0C0F5D5F0C0;
defparam \cp_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \cp_ready~1 (
	.dataa(!in_ready_hold),
	.datab(!in_data_reg_60),
	.datac(!in_narrow_reg),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_ready~1 .extended_lut = "off";
defparam \cp_ready~1 .lut_mask = 64'hC0C0D5C0C0C0D5C0;
defparam \cp_ready~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_burst_uncompressor_5 (
	empty,
	mem_57_0,
	mem_used_0,
	last_packet_beat,
	mem_69_0,
	mem_68_0,
	mem_67_0,
	mem_66_0,
	mem_65_0,
	last_packet_beat1,
	reset,
	last_packet_beat2,
	read,
	clk)/* synthesis synthesis_greybox=0 */;
input 	empty;
input 	mem_57_0;
input 	mem_used_0;
output 	last_packet_beat;
input 	mem_69_0;
input 	mem_68_0;
input 	mem_67_0;
input 	mem_66_0;
input 	mem_65_0;
output 	last_packet_beat1;
input 	reset;
output 	last_packet_beat2;
input 	read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \burst_uncompress_busy~q ;
wire \burst_uncompress_byte_counter~5_combout ;
wire \burst_uncompress_byte_counter[2]~q ;
wire \burst_uncompress_byte_counter~4_combout ;
wire \burst_uncompress_byte_counter[3]~q ;
wire \Add0~2_combout ;
wire \burst_uncompress_byte_counter~3_combout ;
wire \burst_uncompress_byte_counter[4]~q ;
wire \last_packet_beat~3_combout ;
wire \Add1~0_combout ;
wire \burst_uncompress_byte_counter~6_combout ;
wire \burst_uncompress_byte_counter[7]~q ;
wire \burst_uncompress_byte_counter~0_combout ;
wire \Add0~1_combout ;
wire \Add1~1_combout ;
wire \burst_uncompress_byte_counter~2_combout ;
wire \burst_uncompress_byte_counter[5]~q ;
wire \Add0~0_combout ;
wire \burst_uncompress_byte_counter~1_combout ;
wire \burst_uncompress_byte_counter[6]~q ;


cyclonev_lcell_comb \last_packet_beat~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!\burst_uncompress_byte_counter[5]~q ),
	.datad(!\burst_uncompress_byte_counter[4]~q ),
	.datae(!\burst_uncompress_byte_counter[3]~q ),
	.dataf(!\burst_uncompress_byte_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~0 .extended_lut = "off";
defparam \last_packet_beat~0 .lut_mask = 64'h0000000040000000;
defparam \last_packet_beat~0 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~1 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_69_0),
	.datac(!mem_68_0),
	.datad(!mem_67_0),
	.datae(!mem_66_0),
	.dataf(!mem_65_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat1),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~1 .extended_lut = "off";
defparam \last_packet_beat~1 .lut_mask = 64'h0000000080000000;
defparam \last_packet_beat~1 .shared_arith = "off";

cyclonev_lcell_comb \last_packet_beat~2 (
	.dataa(!empty),
	.datab(!mem_57_0),
	.datac(!mem_used_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_packet_beat2),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~2 .extended_lut = "off";
defparam \last_packet_beat~2 .lut_mask = 64'h3331313133313131;
defparam \last_packet_beat~2 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!mem_used_0),
	.datab(!read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h1111111111111111;
defparam \always0~0 .shared_arith = "off";

dffeas burst_uncompress_busy(
	.clk(clk),
	.d(last_packet_beat2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_busy~q ),
	.prn(vcc));
defparam burst_uncompress_busy.is_wysiwyg = "true";
defparam burst_uncompress_busy.power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~5 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~5 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~5 .lut_mask = 64'h00C800FA00C800FA;
defparam \burst_uncompress_byte_counter~5 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[2] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[2]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[2] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[2] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~4 (
	.dataa(!mem_66_0),
	.datab(!mem_65_0),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(!last_packet_beat2),
	.dataf(!\burst_uncompress_byte_counter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~4 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~4 .lut_mask = 64'h000099990000F00F;
defparam \burst_uncompress_byte_counter~4 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[3] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[3]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[3] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\burst_uncompress_byte_counter[4]~q ),
	.datab(!\burst_uncompress_byte_counter[3]~q ),
	.datac(!\burst_uncompress_byte_counter[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6A6A6A6A6A6A6A6A;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~3 (
	.dataa(!mem_67_0),
	.datab(!mem_66_0),
	.datac(!mem_65_0),
	.datad(!last_packet_beat2),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~3 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~3 .lut_mask = 64'h009500FF00950000;
defparam \burst_uncompress_byte_counter~3 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[4] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[4]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[4] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[4] .power_up = "low";

cyclonev_lcell_comb \last_packet_beat~3 (
	.dataa(!\burst_uncompress_byte_counter[6]~q ),
	.datab(!\burst_uncompress_byte_counter[5]~q ),
	.datac(!\burst_uncompress_byte_counter[4]~q ),
	.datad(!\burst_uncompress_byte_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_packet_beat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_packet_beat~3 .extended_lut = "off";
defparam \last_packet_beat~3 .lut_mask = 64'h8000800080008000;
defparam \last_packet_beat~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h8000800080008000;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~6 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~6 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~6 .lut_mask = 64'h0000000C0A0A000C;
defparam \burst_uncompress_byte_counter~6 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[7] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[7]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[7] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[7] .power_up = "low";

cyclonev_lcell_comb \burst_uncompress_byte_counter~0 (
	.dataa(!\burst_uncompress_busy~q ),
	.datab(!\burst_uncompress_byte_counter[2]~q ),
	.datac(!\last_packet_beat~3_combout ),
	.datad(!\burst_uncompress_byte_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~0 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~0 .lut_mask = 64'h5155515551555155;
defparam \burst_uncompress_byte_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!mem_68_0),
	.datab(!mem_67_0),
	.datac(!mem_66_0),
	.datad(!mem_65_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6AAA6AAA6AAA6AAA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~2 (
	.dataa(!last_packet_beat2),
	.datab(!\burst_uncompress_byte_counter~0_combout ),
	.datac(!\Add0~1_combout ),
	.datad(!\Add1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~2 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~2 .lut_mask = 64'h5410541054105410;
defparam \burst_uncompress_byte_counter~2 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[5] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[5]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[5] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\burst_uncompress_byte_counter[5]~q ),
	.datab(!\burst_uncompress_byte_counter[4]~q ),
	.datac(!\burst_uncompress_byte_counter[3]~q ),
	.datad(!\burst_uncompress_byte_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h8000800080008000;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \burst_uncompress_byte_counter~1 (
	.dataa(!mem_69_0),
	.datab(!\burst_uncompress_byte_counter[6]~q ),
	.datac(!last_packet_beat2),
	.datad(!\Add0~0_combout ),
	.datae(!\burst_uncompress_byte_counter~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_uncompress_byte_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_uncompress_byte_counter~1 .extended_lut = "off";
defparam \burst_uncompress_byte_counter~1 .lut_mask = 64'h0505030C0A0A030C;
defparam \burst_uncompress_byte_counter~1 .shared_arith = "off";

dffeas \burst_uncompress_byte_counter[6] (
	.clk(clk),
	.d(\burst_uncompress_byte_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.q(\burst_uncompress_byte_counter[6]~q ),
	.prn(vcc));
defparam \burst_uncompress_byte_counter[6] .is_wysiwyg = "true";
defparam \burst_uncompress_byte_counter[6] .power_up = "low";

endmodule

module terminal_qsys_altera_merlin_slave_translator (
	out_valid_reg,
	in_ready_hold,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	reset,
	m0_write,
	in_data_reg_60,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	out_valid_reg;
input 	in_ready_hold;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	reset;
input 	m0_write;
input 	in_data_reg_60;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h0000044000000440;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_slave_translator_1 (
	in_ready_hold,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	reset,
	m0_write,
	in_data_reg_60,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	reset;
input 	m0_write;
input 	in_data_reg_60;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h0000044000000440;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_slave_translator_2 (
	in_ready_hold,
	out_valid_reg,
	mem_used_1,
	WideOr0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	reset,
	m0_write,
	in_data_reg_60,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	out_valid_reg;
input 	mem_used_1;
input 	WideOr0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
input 	reset;
input 	m0_write;
input 	in_data_reg_60;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;
wire \wait_latency_counter[0]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!WideOr0),
	.datac(!out_valid_reg),
	.datad(!in_data_reg_60),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h0002000200020002;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter[0]~0 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[0]~0 .extended_lut = "off";
defparam \wait_latency_counter[0]~0 .lut_mask = 64'h0015511500155115;
defparam \wait_latency_counter[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0606060606060606;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'h2222222222222222;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!in_ready_hold),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(!\read_latency_shift_reg~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h0000044000000440;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_slave_translator_3 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_30,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_30;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_slave_translator_4 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	av_readdata_pre_10,
	av_readdata_pre_11,
	av_readdata_pre_12,
	av_readdata_pre_13,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_16,
	av_readdata_pre_17,
	av_readdata_pre_18,
	av_readdata_pre_19,
	av_readdata_pre_20,
	av_readdata_pre_21,
	av_readdata_pre_22,
	av_readdata_pre_23,
	av_readdata_pre_24,
	av_readdata_pre_25,
	av_readdata_pre_26,
	av_readdata_pre_27,
	av_readdata_pre_28,
	av_readdata_pre_29,
	av_readdata_pre_30,
	av_readdata_pre_31,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
output 	av_readdata_pre_10;
output 	av_readdata_pre_11;
output 	av_readdata_pre_12;
output 	av_readdata_pre_13;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_16;
output 	av_readdata_pre_17;
output 	av_readdata_pre_18;
output 	av_readdata_pre_19;
output 	av_readdata_pre_20;
output 	av_readdata_pre_21;
output 	av_readdata_pre_22;
output 	av_readdata_pre_23;
output 	av_readdata_pre_24;
output 	av_readdata_pre_25;
output 	av_readdata_pre_26;
output 	av_readdata_pre_27;
output 	av_readdata_pre_28;
output 	av_readdata_pre_29;
output 	av_readdata_pre_30;
output 	av_readdata_pre_31;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_slave_translator_5 (
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_readdata_pre_0,
	av_readdata_pre_1,
	av_readdata_pre_2,
	av_readdata_pre_3,
	av_readdata_pre_4,
	av_readdata_pre_5,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_8,
	av_readdata_pre_9,
	reset,
	write,
	write1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=0 */;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_readdata_pre_0;
output 	av_readdata_pre_1;
output 	av_readdata_pre_2;
output 	av_readdata_pre_3;
output 	av_readdata_pre_4;
output 	av_readdata_pre_5;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_8;
output 	av_readdata_pre_9;
input 	reset;
input 	write;
input 	write1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h0404040404040404;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(gnd),
	.datab(!wait_latency_counter_0),
	.datac(!write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h0C0C0C0C0C0C0C0C;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_traffic_limiter (
	h2f_lw_ARVALID_0,
	h2f_lw_RREADY_0,
	h2f_lw_ARADDR_16,
	h2f_lw_ARADDR_17,
	h2f_lw_ARADDR_18,
	Equal1,
	Equal11,
	cmd_sink_channel,
	sink_ready,
	has_pending_responses1,
	cmd_sink_data,
	sink_ready1,
	WideOr0,
	sink_ready2,
	sink_ready3,
	cmd_sink_ready,
	src_payload_0,
	WideOr1,
	last_channel_5,
	WideOr01,
	reset,
	last_channel_3,
	last_channel_0,
	last_channel_1,
	last_channel_2,
	last_channel_4,
	WideOr02,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_RREADY_0;
input 	h2f_lw_ARADDR_16;
input 	h2f_lw_ARADDR_17;
input 	h2f_lw_ARADDR_18;
input 	Equal1;
input 	Equal11;
input 	[5:0] cmd_sink_channel;
input 	sink_ready;
output 	has_pending_responses1;
input 	[115:0] cmd_sink_data;
input 	sink_ready1;
input 	WideOr0;
input 	sink_ready2;
input 	sink_ready3;
output 	cmd_sink_ready;
input 	src_payload_0;
input 	WideOr1;
output 	last_channel_5;
input 	WideOr01;
input 	reset;
output 	last_channel_3;
output 	last_channel_0;
output 	last_channel_1;
output 	last_channel_2;
output 	last_channel_4;
input 	WideOr02;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~combout ;
wire \last_dest_id[0]~q ;
wire \last_dest_id[1]~q ;
wire \Equal0~0_combout ;
wire \last_dest_id[2]~q ;
wire \Equal0~1_combout ;
wire \internal_valid~1_combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \internal_valid~0_combout ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

cyclonev_lcell_comb \cmd_sink_ready~0 (
	.dataa(!sink_ready),
	.datab(!\internal_valid~0_combout ),
	.datac(!sink_ready1),
	.datad(!WideOr0),
	.datae(!sink_ready2),
	.dataf(!sink_ready3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cmd_sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_sink_ready~0 .extended_lut = "off";
defparam \cmd_sink_ready~0 .lut_mask = 64'hCC4CCCCCCCCCCCCC;
defparam \cmd_sink_ready~0 .shared_arith = "off";

dffeas \last_channel[5] (
	.clk(clk),
	.d(cmd_sink_channel[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(last_channel_5),
	.prn(vcc));
defparam \last_channel[5] .is_wysiwyg = "true";
defparam \last_channel[5] .power_up = "low";

dffeas \last_channel[3] (
	.clk(clk),
	.d(cmd_sink_channel[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(last_channel_3),
	.prn(vcc));
defparam \last_channel[3] .is_wysiwyg = "true";
defparam \last_channel[3] .power_up = "low";

dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas \last_channel[1] (
	.clk(clk),
	.d(cmd_sink_channel[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(last_channel_1),
	.prn(vcc));
defparam \last_channel[1] .is_wysiwyg = "true";
defparam \last_channel[1] .power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

dffeas \last_channel[4] (
	.clk(clk),
	.d(cmd_sink_channel[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(last_channel_4),
	.prn(vcc));
defparam \last_channel[4] .is_wysiwyg = "true";
defparam \last_channel[4] .power_up = "low";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb response_sink_accepted(
	.dataa(!h2f_lw_RREADY_0),
	.datab(!src_payload_0),
	.datac(!WideOr1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam response_sink_accepted.extended_lut = "off";
defparam response_sink_accepted.lut_mask = 64'h0101010101010101;
defparam response_sink_accepted.shared_arith = "off";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[89]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(\last_dest_id[0]~q ),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(cmd_sink_data[90]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(\last_dest_id[1]~q ),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!h2f_lw_ARADDR_18),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(!\last_dest_id[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFC50000003A;
defparam \Equal0~0 .shared_arith = "off";

dffeas \last_dest_id[2] (
	.clk(clk),
	.d(cmd_sink_data[91]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~1_combout ),
	.q(\last_dest_id[2]~q ),
	.prn(vcc));
defparam \last_dest_id[2] .is_wysiwyg = "true";
defparam \last_dest_id[2] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(gnd),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(!\last_dest_id[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h00000022FFFFFFDD;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \internal_valid~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses1),
	.datac(!\last_dest_id[0]~q ),
	.datad(!cmd_sink_data[89]),
	.datae(!\Equal0~0_combout ),
	.dataf(!\Equal0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_valid~1 .extended_lut = "off";
defparam \internal_valid~1 .lut_mask = 64'h5445444444444444;
defparam \internal_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!sink_ready1),
	.datab(!WideOr02),
	.datac(!sink_ready2),
	.datad(!sink_ready3),
	.datae(!\response_sink_accepted~combout ),
	.dataf(!\internal_valid~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h0000FFFFDFFF2000;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[1]~q ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6969696969696969;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!WideOr01),
	.datac(!\pending_response_count[1]~q ),
	.datad(!\pending_response_count[0]~q ),
	.datae(!\response_sink_accepted~combout ),
	.dataf(!\internal_valid~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h55555505D5555545;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \internal_valid~0 (
	.dataa(!has_pending_responses1),
	.datab(!\last_dest_id[0]~q ),
	.datac(!cmd_sink_data[89]),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_valid~0 .extended_lut = "off";
defparam \internal_valid~0 .lut_mask = 64'h1455555514555555;
defparam \internal_valid~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_traffic_limiter_1 (
	h2f_lw_BREADY_0,
	h2f_lw_WLAST_0,
	write_addr_data_both_valid,
	Equal3,
	Equal31,
	Equal4,
	has_pending_responses1,
	last_channel_2,
	last_channel_4,
	sink_ready,
	sink_ready1,
	sink_ready2,
	nonposted_cmd_accepted,
	src0_valid,
	mem_57_0,
	src0_valid1,
	mem_57_01,
	src0_valid2,
	WideOr1,
	comb,
	mem_117_0,
	last_packet_beat,
	last_packet_beat1,
	comb1,
	mem_117_01,
	last_packet_beat2,
	last_packet_beat3,
	nonposted_cmd_accepted1,
	reset,
	last_channel_3,
	cmd_sink_channel,
	WideOr0,
	src_payload,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_WLAST_0;
input 	write_addr_data_both_valid;
input 	Equal3;
input 	Equal31;
input 	Equal4;
output 	has_pending_responses1;
output 	last_channel_2;
output 	last_channel_4;
input 	sink_ready;
input 	sink_ready1;
input 	sink_ready2;
output 	nonposted_cmd_accepted;
input 	src0_valid;
input 	mem_57_0;
input 	src0_valid1;
input 	mem_57_01;
input 	src0_valid2;
input 	WideOr1;
input 	comb;
input 	mem_117_0;
input 	last_packet_beat;
input 	last_packet_beat1;
input 	comb1;
input 	mem_117_01;
input 	last_packet_beat2;
input 	last_packet_beat3;
output 	nonposted_cmd_accepted1;
input 	reset;
output 	last_channel_3;
input 	[5:0] cmd_sink_channel;
input 	WideOr0;
input 	src_payload;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \suppress_change_dest_id~0_combout ;
wire \internal_valid~0_combout ;
wire \pending_response_count[0]~1_combout ;
wire \response_sink_accepted~0_combout ;
wire \response_sink_accepted~1_combout ;
wire \response_sink_accepted~2_combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~1_combout ;
wire \has_pending_responses~2_combout ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~0_combout ),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

dffeas \last_channel[4] (
	.clk(clk),
	.d(cmd_sink_channel[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~0_combout ),
	.q(last_channel_4),
	.prn(vcc));
defparam \last_channel[4] .is_wysiwyg = "true";
defparam \last_channel[4] .power_up = "low";

cyclonev_lcell_comb \nonposted_cmd_accepted~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!write_addr_data_both_valid),
	.datac(!\suppress_change_dest_id~0_combout ),
	.datad(!sink_ready),
	.datae(!sink_ready1),
	.dataf(!sink_ready2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted),
	.sumout(),
	.cout(),
	.shareout());
defparam \nonposted_cmd_accepted~0 .extended_lut = "off";
defparam \nonposted_cmd_accepted~0 .lut_mask = 64'h0010101010101010;
defparam \nonposted_cmd_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \nonposted_cmd_accepted~1 (
	.dataa(!write_addr_data_both_valid),
	.datab(!\suppress_change_dest_id~0_combout ),
	.datac(!sink_ready),
	.datad(!sink_ready1),
	.datae(!sink_ready2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam \nonposted_cmd_accepted~1 .extended_lut = "off";
defparam \nonposted_cmd_accepted~1 .lut_mask = 64'h0444444404444444;
defparam \nonposted_cmd_accepted~1 .shared_arith = "off";

dffeas \last_channel[3] (
	.clk(clk),
	.d(cmd_sink_channel[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_valid~0_combout ),
	.q(last_channel_3),
	.prn(vcc));
defparam \last_channel[3] .is_wysiwyg = "true";
defparam \last_channel[3] .power_up = "low";

cyclonev_lcell_comb \suppress_change_dest_id~0 (
	.dataa(!Equal3),
	.datab(!Equal31),
	.datac(!Equal4),
	.datad(!has_pending_responses1),
	.datae(!last_channel_2),
	.dataf(!last_channel_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\suppress_change_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~0 .extended_lut = "off";
defparam \suppress_change_dest_id~0 .lut_mask = 64'h00FB00EE001500FF;
defparam \suppress_change_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \internal_valid~0 (
	.dataa(!write_addr_data_both_valid),
	.datab(!\suppress_change_dest_id~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_valid~0 .extended_lut = "off";
defparam \internal_valid~0 .lut_mask = 64'h4444444444444444;
defparam \internal_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~1 (
	.dataa(!\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~1 .extended_lut = "off";
defparam \pending_response_count[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \pending_response_count[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!src0_valid1),
	.datad(!mem_117_0),
	.datae(!last_packet_beat),
	.dataf(!last_packet_beat1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h000C000D000D000D;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~1 (
	.dataa(!comb1),
	.datab(!mem_57_01),
	.datac(!src0_valid2),
	.datad(!mem_117_01),
	.datae(!last_packet_beat2),
	.dataf(!last_packet_beat3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~1 .extended_lut = "off";
defparam \response_sink_accepted~1 .lut_mask = 64'h000C000D000D000D;
defparam \response_sink_accepted~1 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~2 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!src0_valid),
	.datac(!src_payload),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(!\response_sink_accepted~1_combout ),
	.dataf(!WideOr1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~2 .extended_lut = "off";
defparam \response_sink_accepted~2 .lut_mask = 64'h0000000001555555;
defparam \response_sink_accepted~2 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[1]~0 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!\internal_valid~0_combout ),
	.datac(!sink_ready),
	.datad(!WideOr0),
	.datae(!\response_sink_accepted~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[1]~0 .extended_lut = "off";
defparam \pending_response_count[1]~0 .lut_mask = 64'h1101EEFE1101EEFE;
defparam \pending_response_count[1]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\pending_response_count[1]~q ),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6969696969696969;
defparam \Add0~0 .shared_arith = "off";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!\pending_response_count[1]~q ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'h5551555155515551;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~1 (
	.dataa(!has_pending_responses1),
	.datab(!\pending_response_count[1]~q ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~1 .extended_lut = "off";
defparam \has_pending_responses~1 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \has_pending_responses~1 .shared_arith = "off";

cyclonev_lcell_comb \has_pending_responses~2 (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!\internal_valid~0_combout ),
	.datac(!sink_ready),
	.datad(!WideOr0),
	.datae(!\has_pending_responses~0_combout ),
	.dataf(!\has_pending_responses~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~2 .extended_lut = "off";
defparam \has_pending_responses~2 .lut_mask = 64'h1101FFFF0000FFFF;
defparam \has_pending_responses~2 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_demux (
	h2f_lw_AWVALID_0,
	h2f_lw_WVALID_0,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	nxt_in_ready3,
	nxt_in_ready4,
	nxt_in_ready5,
	Equal3,
	Equal31,
	Equal4,
	has_pending_responses,
	last_channel_2,
	last_channel_4,
	saved_grant_0,
	sink_ready,
	saved_grant_01,
	sink_ready1,
	saved_grant_02,
	sink_ready2,
	last_channel_3,
	src3_valid,
	src2_valid,
	src4_valid,
	src4_valid1,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWVALID_0;
input 	h2f_lw_WVALID_0;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	nxt_in_ready3;
input 	nxt_in_ready4;
input 	nxt_in_ready5;
input 	Equal3;
input 	Equal31;
input 	Equal4;
input 	has_pending_responses;
input 	last_channel_2;
input 	last_channel_4;
input 	saved_grant_0;
output 	sink_ready;
input 	saved_grant_01;
output 	sink_ready1;
input 	saved_grant_02;
output 	sink_ready2;
input 	last_channel_3;
output 	src3_valid;
output 	src2_valid;
output 	src4_valid;
output 	src4_valid1;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~3_combout ;
wire \sink_ready~4_combout ;


cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!nxt_in_ready3),
	.datab(!nxt_in_ready2),
	.datac(!saved_grant_0),
	.datad(!Equal3),
	.datae(!Equal4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h0000000700000007;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!nxt_in_ready4),
	.datab(!nxt_in_ready1),
	.datac(!saved_grant_01),
	.datad(!Equal3),
	.datae(!Equal31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'h0000000700000007;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!nxt_in_ready5),
	.datab(!nxt_in_ready),
	.datac(!saved_grant_02),
	.datad(!Equal3),
	.datae(!Equal31),
	.dataf(!Equal4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'h0707070007000700;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \src3_valid~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!has_pending_responses),
	.datad(!last_channel_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src3_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~0 .extended_lut = "off";
defparam \src3_valid~0 .lut_mask = 64'h1011101110111011;
defparam \src3_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!has_pending_responses),
	.datad(!last_channel_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'h1011101110111011;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src4_valid~0 (
	.dataa(!Equal3),
	.datab(!Equal31),
	.datac(!Equal4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src4_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src4_valid~0 .extended_lut = "off";
defparam \src4_valid~0 .lut_mask = 64'hEAEAEAEAEAEAEAEA;
defparam \src4_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src4_valid~1 (
	.dataa(!h2f_lw_AWVALID_0),
	.datab(!h2f_lw_WVALID_0),
	.datac(!has_pending_responses),
	.datad(!last_channel_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src4_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src4_valid~1 .extended_lut = "off";
defparam \src4_valid~1 .lut_mask = 64'h1011101110111011;
defparam \src4_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!nxt_in_ready4),
	.datab(!nxt_in_ready1),
	.datac(!nxt_in_ready5),
	.datad(!nxt_in_ready),
	.datae(!\sink_ready~3_combout ),
	.dataf(!\sink_ready~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hFFFF8888F0008000;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!saved_grant_01),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'h0101010101010101;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!saved_grant_02),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(!Equal4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'h5444544454445444;
defparam \sink_ready~4 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_demux_1 (
	h2f_lw_ARVALID_0,
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_16,
	h2f_lw_ARADDR_17,
	h2f_lw_ARADDR_18,
	nxt_in_ready,
	nxt_in_ready1,
	nxt_in_ready2,
	Equal1,
	Equal11,
	Equal5,
	saved_grant_1,
	nxt_in_ready3,
	nxt_in_ready4,
	sink_ready,
	has_pending_responses,
	saved_grant_11,
	Equal4,
	Equal41,
	nxt_in_ready5,
	sink_ready1,
	nxt_in_ready6,
	nxt_in_ready7,
	saved_grant_12,
	Equal12,
	nxt_in_ready8,
	nxt_in_ready9,
	saved_grant_13,
	WideOr01,
	saved_grant_14,
	Equal3,
	nxt_in_ready10,
	sink_ready2,
	saved_grant_15,
	nxt_in_ready11,
	src_channel_4,
	sink_ready3,
	WideOr02,
	last_channel_3,
	src3_valid,
	src3_valid1,
	last_channel_2,
	src2_valid,
	src2_valid1,
	last_channel_4,
	src4_valid,
	WideOr03,
	src4_valid1)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_16;
input 	h2f_lw_ARADDR_17;
input 	h2f_lw_ARADDR_18;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	nxt_in_ready2;
input 	Equal1;
input 	Equal11;
input 	Equal5;
input 	saved_grant_1;
input 	nxt_in_ready3;
input 	nxt_in_ready4;
output 	sink_ready;
input 	has_pending_responses;
input 	saved_grant_11;
input 	Equal4;
input 	Equal41;
input 	nxt_in_ready5;
output 	sink_ready1;
input 	nxt_in_ready6;
input 	nxt_in_ready7;
input 	saved_grant_12;
input 	Equal12;
input 	nxt_in_ready8;
input 	nxt_in_ready9;
input 	saved_grant_13;
output 	WideOr01;
input 	saved_grant_14;
input 	Equal3;
input 	nxt_in_ready10;
output 	sink_ready2;
input 	saved_grant_15;
input 	nxt_in_ready11;
input 	src_channel_4;
output 	sink_ready3;
output 	WideOr02;
input 	last_channel_3;
output 	src3_valid;
output 	src3_valid1;
input 	last_channel_2;
output 	src2_valid;
output 	src2_valid1;
input 	last_channel_4;
output 	src4_valid;
output 	WideOr03;
output 	src4_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~2_combout ;
wire \sink_ready~3_combout ;


cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!Equal5),
	.datab(!saved_grant_1),
	.datac(!nxt_in_ready3),
	.datad(!nxt_in_ready4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'h1101110111011101;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!saved_grant_11),
	.datab(!Equal41),
	.datac(!nxt_in_ready5),
	.datad(!nxt_in_ready2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'h0111011101110111;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!nxt_in_ready6),
	.datab(!nxt_in_ready7),
	.datac(!\sink_ready~2_combout ),
	.datad(!nxt_in_ready8),
	.datae(!nxt_in_ready9),
	.dataf(!\sink_ready~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF2F2F2F20000F200;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!saved_grant_14),
	.datab(!Equal3),
	.datac(!nxt_in_ready10),
	.datad(!nxt_in_ready1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'h0111011101110111;
defparam \sink_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~5 (
	.dataa(!saved_grant_15),
	.datab(!nxt_in_ready11),
	.datac(!nxt_in_ready),
	.datad(!src_channel_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~5 .extended_lut = "off";
defparam \sink_ready~5 .lut_mask = 64'h0015001500150015;
defparam \sink_ready~5 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!sink_ready),
	.datab(!sink_ready1),
	.datac(!WideOr01),
	.datad(!sink_ready2),
	.datae(!sink_ready3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr02),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h0800000008000000;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \src3_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src3_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~0 .extended_lut = "off";
defparam \src3_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src3_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src3_valid~1 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!Equal4),
	.datae(!src3_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src3_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~1 .extended_lut = "off";
defparam \src3_valid~1 .lut_mask = 64'h0000000200000002;
defparam \src3_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~1 (
	.dataa(!h2f_lw_ARADDR_17),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!Equal12),
	.datae(!src2_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~1 .extended_lut = "off";
defparam \src2_valid~1 .lut_mask = 64'h0000000100000001;
defparam \src2_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src4_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!src_channel_4),
	.datad(!last_channel_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src4_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src4_valid~0 .extended_lut = "off";
defparam \src4_valid~0 .lut_mask = 64'h0405040504050405;
defparam \src4_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!sink_ready),
	.datab(!WideOr01),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr03),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'h2222222222222222;
defparam \WideOr0~1 .shared_arith = "off";

cyclonev_lcell_comb \src4_valid~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src4_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src4_valid~1 .extended_lut = "off";
defparam \src4_valid~1 .lut_mask = 64'h4545454545454545;
defparam \src4_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!saved_grant_12),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(!Equal12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'h0000000000000008;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!h2f_lw_ARADDR_18),
	.datad(!saved_grant_13),
	.datae(!Equal1),
	.dataf(!Equal11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'h0000000000000020;
defparam \sink_ready~3 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux (
	h2f_lw_ARVALID_0,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	has_pending_responses,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Equal1,
	last_channel_0,
	src_valid,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	has_pending_responses;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal1;
input 	last_channel_0;
output 	src_valid;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h4545454545454545;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!saved_grant_1),
	.datab(!Equal1),
	.datac(!nxt_in_ready),
	.datad(!nxt_in_ready1),
	.datae(!\packet_in_progress~q ),
	.dataf(!src_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h0000FFFF0010EEFE;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!saved_grant_1),
	.datab(!Equal1),
	.datac(!\packet_in_progress~q ),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h0535053505350535;
defparam \saved_grant[1]~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_1 (
	h2f_lw_ARVALID_0,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	has_pending_responses,
	nxt_in_ready,
	nxt_in_ready1,
	saved_grant_1,
	altera_reset_synchronizer_int_chain_out,
	Equal2,
	last_channel_1,
	src_valid,
	src_valid1,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	has_pending_responses;
input 	nxt_in_ready;
input 	nxt_in_ready1;
output 	saved_grant_1;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal2;
input 	last_channel_1;
output 	src_valid;
output 	src_valid1;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~0_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!saved_grant_1),
	.datac(!Equal2),
	.datad(!has_pending_responses),
	.datae(!last_channel_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0100010101000101;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h4545454545454545;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!nxt_in_ready),
	.datab(!nxt_in_ready1),
	.datac(!\packet_in_progress~q ),
	.datad(!src_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h0F220F220F220F22;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!saved_grant_1),
	.datab(!Equal2),
	.datac(!\packet_in_progress~q ),
	.datad(!src_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h0535053505350535;
defparam \saved_grant[1]~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_2 (
	h2f_lw_WLAST_0,
	h2f_lw_ARADDR_17,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	nxt_in_ready,
	Equal1,
	Equal11,
	Equal12,
	saved_grant_1,
	nxt_in_ready1,
	Equal3,
	Equal31,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	src2_valid,
	src2_valid1,
	src2_valid2,
	src_valid,
	src_payload_0,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_73,
	src_data_72,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	src_data_77,
	Selector5,
	Selector12,
	src_data_71,
	Selector6,
	nxt_out_burstwrap_0,
	src_data_70,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_ARADDR_17;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	nxt_in_ready;
input 	Equal1;
input 	Equal11;
input 	Equal12;
output 	saved_grant_1;
input 	nxt_in_ready1;
input 	Equal3;
input 	Equal31;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src2_valid;
input 	src2_valid1;
input 	src2_valid2;
output 	src_valid;
output 	src_payload_0;
output 	src_data_78;
output 	src_data_79;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_73;
output 	src_data_72;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_100;
output 	src_data_101;
output 	src_data_102;
output 	src_data_103;
output 	src_data_77;
input 	Selector5;
input 	Selector12;
output 	src_data_71;
input 	Selector6;
input 	nxt_out_burstwrap_0;
output 	src_data_70;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


terminal_qsys_altera_merlin_arbitrator_1 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal3(Equal3),
	.Equal31(Equal31),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src2_valid(src2_valid),
	.src2_valid1(src2_valid2),
	.grant_1(\arb|grant[1]~0_combout ),
	.WideOr1(\WideOr1~combout ),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_ARADDR_17),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!saved_grant_1),
	.datae(!Equal12),
	.dataf(!src2_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0000000000000001;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73] .extended_lut = "off";
defparam \src_data[73] .lut_mask = 64'h3075307530753075;
defparam \src_data[73] .shared_arith = "off";

cyclonev_lcell_comb \src_data[72] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72] .extended_lut = "off";
defparam \src_data[72] .lut_mask = 64'h3075307530753075;
defparam \src_data[72] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_WDATA_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_WDATA_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!h2f_lw_WDATA_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!h2f_lw_WDATA_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!h2f_lw_WDATA_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!h2f_lw_WDATA_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!h2f_lw_WDATA_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!h2f_lw_WDATA_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!h2f_lw_WDATA_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!h2f_lw_WDATA_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!h2f_lw_WDATA_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!h2f_lw_WDATA_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!h2f_lw_WDATA_28),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!h2f_lw_WDATA_29),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!h2f_lw_WDATA_30),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h1111111111111111;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!h2f_lw_WDATA_31),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[100] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_100),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100] .extended_lut = "off";
defparam \src_data[100] .lut_mask = 64'h0537053705370537;
defparam \src_data[100] .shared_arith = "off";

cyclonev_lcell_comb \src_data[101] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101] .extended_lut = "off";
defparam \src_data[101] .lut_mask = 64'h0537053705370537;
defparam \src_data[101] .shared_arith = "off";

cyclonev_lcell_comb \src_data[102] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102] .extended_lut = "off";
defparam \src_data[102] .lut_mask = 64'h0537053705370537;
defparam \src_data[102] .shared_arith = "off";

cyclonev_lcell_comb \src_data[103] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103] .extended_lut = "off";
defparam \src_data[103] .lut_mask = 64'h0537053705370537;
defparam \src_data[103] .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_data[71] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71] .extended_lut = "off";
defparam \src_data[71] .lut_mask = 64'h3075307530753075;
defparam \src_data[71] .shared_arith = "off";

cyclonev_lcell_comb \src_data[70] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!nxt_out_burstwrap_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70] .extended_lut = "off";
defparam \src_data[70] .lut_mask = 64'h3075307530753075;
defparam \src_data[70] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_0),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(!src2_valid),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!\WideOr1~combout ),
	.datad(!src_payload_0),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'h0F7F00700F7F0070;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_arbitrator_1 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal3,
	Equal31,
	reset,
	src2_valid,
	src2_valid1,
	grant_1,
	WideOr1,
	src_payload_0,
	packet_in_progress,
	grant_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal3;
input 	Equal31;
input 	reset;
input 	src2_valid;
input 	src2_valid1;
output 	grant_1;
input 	WideOr1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!Equal3),
	.datab(!Equal31),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!src2_valid),
	.dataf(!src2_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00000000FF0FEF0F;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!Equal3),
	.datab(!Equal31),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!src2_valid),
	.dataf(!src2_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0000110100001100;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal3),
	.datab(!Equal31),
	.datac(!src2_valid),
	.datad(!src2_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_3 (
	h2f_lw_WLAST_0,
	h2f_lw_ARADDR_16,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WDATA_10,
	h2f_lw_WDATA_11,
	h2f_lw_WDATA_12,
	h2f_lw_WDATA_13,
	h2f_lw_WDATA_14,
	h2f_lw_WDATA_15,
	h2f_lw_WDATA_16,
	h2f_lw_WDATA_17,
	h2f_lw_WDATA_18,
	h2f_lw_WDATA_19,
	h2f_lw_WDATA_20,
	h2f_lw_WDATA_21,
	h2f_lw_WDATA_22,
	h2f_lw_WDATA_23,
	h2f_lw_WDATA_24,
	h2f_lw_WDATA_25,
	h2f_lw_WDATA_26,
	h2f_lw_WDATA_27,
	h2f_lw_WDATA_28,
	h2f_lw_WDATA_29,
	h2f_lw_WDATA_30,
	h2f_lw_WDATA_31,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	nxt_in_ready,
	Equal1,
	Equal11,
	saved_grant_1,
	Equal4,
	nxt_in_ready1,
	Equal3,
	Equal41,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	src3_valid,
	src3_valid1,
	src3_valid2,
	src_valid,
	src_payload_0,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	src_payload,
	Selector3,
	Selector10,
	src_data_73,
	Selector4,
	Selector11,
	src_data_72,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	src_data_77,
	Selector5,
	Selector12,
	src_data_71,
	Selector6,
	nxt_out_burstwrap_0,
	src_data_70,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_ARADDR_16;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WDATA_10;
input 	h2f_lw_WDATA_11;
input 	h2f_lw_WDATA_12;
input 	h2f_lw_WDATA_13;
input 	h2f_lw_WDATA_14;
input 	h2f_lw_WDATA_15;
input 	h2f_lw_WDATA_16;
input 	h2f_lw_WDATA_17;
input 	h2f_lw_WDATA_18;
input 	h2f_lw_WDATA_19;
input 	h2f_lw_WDATA_20;
input 	h2f_lw_WDATA_21;
input 	h2f_lw_WDATA_22;
input 	h2f_lw_WDATA_23;
input 	h2f_lw_WDATA_24;
input 	h2f_lw_WDATA_25;
input 	h2f_lw_WDATA_26;
input 	h2f_lw_WDATA_27;
input 	h2f_lw_WDATA_28;
input 	h2f_lw_WDATA_29;
input 	h2f_lw_WDATA_30;
input 	h2f_lw_WDATA_31;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	nxt_in_ready;
input 	Equal1;
input 	Equal11;
output 	saved_grant_1;
input 	Equal4;
input 	nxt_in_ready1;
input 	Equal3;
input 	Equal41;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src3_valid;
input 	src3_valid1;
input 	src3_valid2;
output 	src_valid;
output 	src_payload_0;
output 	src_data_78;
output 	src_data_79;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
output 	src_payload;
input 	Selector3;
input 	Selector10;
output 	src_data_73;
input 	Selector4;
input 	Selector11;
output 	src_data_72;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_100;
output 	src_data_101;
output 	src_data_102;
output 	src_data_103;
output 	src_data_77;
input 	Selector5;
input 	Selector12;
output 	src_data_71;
input 	Selector6;
input 	nxt_out_burstwrap_0;
output 	src_data_70;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \WideOr1~combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


terminal_qsys_altera_merlin_arbitrator_2 arb(
	.nxt_in_ready(nxt_in_ready),
	.nxt_in_ready1(nxt_in_ready1),
	.Equal3(Equal3),
	.Equal4(Equal41),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src3_valid(src3_valid),
	.src3_valid1(src3_valid2),
	.grant_1(\arb|grant[1]~0_combout ),
	.WideOr1(\WideOr1~combout ),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!saved_grant_1),
	.datae(!Equal4),
	.dataf(!src3_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0000000000000002;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73] .extended_lut = "off";
defparam \src_data[73] .lut_mask = 64'h3075307530753075;
defparam \src_data[73] .shared_arith = "off";

cyclonev_lcell_comb \src_data[72] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72] .extended_lut = "off";
defparam \src_data[72] .lut_mask = 64'h3075307530753075;
defparam \src_data[72] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!h2f_lw_WDATA_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h1111111111111111;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!h2f_lw_WDATA_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h1111111111111111;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!h2f_lw_WDATA_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h1111111111111111;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!h2f_lw_WDATA_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h1111111111111111;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!h2f_lw_WDATA_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h1111111111111111;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!h2f_lw_WDATA_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h1111111111111111;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!h2f_lw_WDATA_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h1111111111111111;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!h2f_lw_WDATA_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h1111111111111111;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!h2f_lw_WDATA_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h1111111111111111;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!h2f_lw_WDATA_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h1111111111111111;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!h2f_lw_WDATA_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h1111111111111111;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!h2f_lw_WDATA_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h1111111111111111;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!h2f_lw_WDATA_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h1111111111111111;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!h2f_lw_WDATA_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h1111111111111111;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!h2f_lw_WDATA_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h1111111111111111;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!h2f_lw_WDATA_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h1111111111111111;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!h2f_lw_WDATA_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h1111111111111111;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!h2f_lw_WDATA_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h1111111111111111;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!h2f_lw_WDATA_28),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h1111111111111111;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!h2f_lw_WDATA_29),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h1111111111111111;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!h2f_lw_WDATA_30),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h1111111111111111;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!h2f_lw_WDATA_31),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h1111111111111111;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[100] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_100),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100] .extended_lut = "off";
defparam \src_data[100] .lut_mask = 64'h0537053705370537;
defparam \src_data[100] .shared_arith = "off";

cyclonev_lcell_comb \src_data[101] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101] .extended_lut = "off";
defparam \src_data[101] .lut_mask = 64'h0537053705370537;
defparam \src_data[101] .shared_arith = "off";

cyclonev_lcell_comb \src_data[102] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102] .extended_lut = "off";
defparam \src_data[102] .lut_mask = 64'h0537053705370537;
defparam \src_data[102] .shared_arith = "off";

cyclonev_lcell_comb \src_data[103] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103] .extended_lut = "off";
defparam \src_data[103] .lut_mask = 64'h0537053705370537;
defparam \src_data[103] .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_data[71] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71] .extended_lut = "off";
defparam \src_data[71] .lut_mask = 64'h3075307530753075;
defparam \src_data[71] .shared_arith = "off";

cyclonev_lcell_comb \src_data[70] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!nxt_out_burstwrap_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70] .extended_lut = "off";
defparam \src_data[70] .lut_mask = 64'h3075307530753075;
defparam \src_data[70] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!saved_grant_0),
	.datab(!Equal3),
	.datac(!Equal41),
	.datad(!src3_valid),
	.datae(!src_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFE0000FFFE0000;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!\WideOr1~combout ),
	.datad(!src_payload_0),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'h0F7F00700F7F0070;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_arbitrator_2 (
	nxt_in_ready,
	nxt_in_ready1,
	Equal3,
	Equal4,
	reset,
	src3_valid,
	src3_valid1,
	grant_1,
	WideOr1,
	src_payload_0,
	packet_in_progress,
	grant_0,
	clk)/* synthesis synthesis_greybox=0 */;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	Equal3;
input 	Equal4;
input 	reset;
input 	src3_valid;
input 	src3_valid1;
output 	grant_1;
input 	WideOr1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!Equal3),
	.datab(!Equal4),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!src3_valid),
	.dataf(!src3_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h00000000FF0FEF0F;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!Equal3),
	.datab(!Equal4),
	.datac(!\top_priority_reg[1]~q ),
	.datad(!\top_priority_reg[0]~q ),
	.datae(!src3_valid),
	.dataf(!src3_valid1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0000110100001100;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!Equal3),
	.datab(!Equal4),
	.datac(!src3_valid),
	.datad(!src3_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!WideOr1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h0F7F007000000000;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_4 (
	h2f_lw_ARVALID_0,
	h2f_lw_WLAST_0,
	h2f_lw_ARID_0,
	h2f_lw_ARID_1,
	h2f_lw_ARID_2,
	h2f_lw_ARID_3,
	h2f_lw_ARID_4,
	h2f_lw_ARID_5,
	h2f_lw_ARID_6,
	h2f_lw_ARID_7,
	h2f_lw_ARID_8,
	h2f_lw_ARID_9,
	h2f_lw_ARID_10,
	h2f_lw_ARID_11,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	h2f_lw_AWID_0,
	h2f_lw_AWID_1,
	h2f_lw_AWID_2,
	h2f_lw_AWID_3,
	h2f_lw_AWID_4,
	h2f_lw_AWID_5,
	h2f_lw_AWID_6,
	h2f_lw_AWID_7,
	h2f_lw_AWID_8,
	h2f_lw_AWID_9,
	h2f_lw_AWID_10,
	h2f_lw_AWID_11,
	h2f_lw_AWSIZE_0,
	h2f_lw_AWSIZE_1,
	h2f_lw_AWSIZE_2,
	h2f_lw_WDATA_0,
	h2f_lw_WDATA_1,
	h2f_lw_WDATA_2,
	h2f_lw_WDATA_3,
	h2f_lw_WDATA_4,
	h2f_lw_WDATA_5,
	h2f_lw_WDATA_6,
	h2f_lw_WDATA_7,
	h2f_lw_WDATA_8,
	h2f_lw_WDATA_9,
	h2f_lw_WSTRB_0,
	h2f_lw_WSTRB_1,
	h2f_lw_WSTRB_2,
	h2f_lw_WSTRB_3,
	nxt_in_ready,
	has_pending_responses,
	saved_grant_1,
	nxt_in_ready1,
	src_channel_4,
	Equal3,
	Equal31,
	Equal4,
	saved_grant_0,
	altera_reset_synchronizer_int_chain_out,
	src4_valid,
	src4_valid1,
	last_channel_4,
	src4_valid2,
	src_valid,
	src_valid1,
	src_payload_0,
	src_data_78,
	src_data_79,
	src_data_35,
	src_data_34,
	src_data_33,
	src_data_32,
	Selector3,
	Selector10,
	Selector4,
	Selector11,
	src_payload,
	src_data_73,
	src_data_72,
	src_payload1,
	src_payload2,
	src_payload3,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	nxt_in_ready2,
	src4_valid3,
	src_data_92,
	src_data_93,
	src_data_94,
	src_data_95,
	src_data_96,
	src_data_97,
	src_data_98,
	src_data_99,
	src_data_100,
	src_data_101,
	src_data_102,
	src_data_103,
	src_data_77,
	Selector5,
	Selector12,
	src_data_71,
	Selector6,
	nxt_out_burstwrap_0,
	src_data_70,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_WLAST_0;
input 	h2f_lw_ARID_0;
input 	h2f_lw_ARID_1;
input 	h2f_lw_ARID_2;
input 	h2f_lw_ARID_3;
input 	h2f_lw_ARID_4;
input 	h2f_lw_ARID_5;
input 	h2f_lw_ARID_6;
input 	h2f_lw_ARID_7;
input 	h2f_lw_ARID_8;
input 	h2f_lw_ARID_9;
input 	h2f_lw_ARID_10;
input 	h2f_lw_ARID_11;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	h2f_lw_AWID_0;
input 	h2f_lw_AWID_1;
input 	h2f_lw_AWID_2;
input 	h2f_lw_AWID_3;
input 	h2f_lw_AWID_4;
input 	h2f_lw_AWID_5;
input 	h2f_lw_AWID_6;
input 	h2f_lw_AWID_7;
input 	h2f_lw_AWID_8;
input 	h2f_lw_AWID_9;
input 	h2f_lw_AWID_10;
input 	h2f_lw_AWID_11;
input 	h2f_lw_AWSIZE_0;
input 	h2f_lw_AWSIZE_1;
input 	h2f_lw_AWSIZE_2;
input 	h2f_lw_WDATA_0;
input 	h2f_lw_WDATA_1;
input 	h2f_lw_WDATA_2;
input 	h2f_lw_WDATA_3;
input 	h2f_lw_WDATA_4;
input 	h2f_lw_WDATA_5;
input 	h2f_lw_WDATA_6;
input 	h2f_lw_WDATA_7;
input 	h2f_lw_WDATA_8;
input 	h2f_lw_WDATA_9;
input 	h2f_lw_WSTRB_0;
input 	h2f_lw_WSTRB_1;
input 	h2f_lw_WSTRB_2;
input 	h2f_lw_WSTRB_3;
input 	nxt_in_ready;
input 	has_pending_responses;
output 	saved_grant_1;
input 	nxt_in_ready1;
input 	src_channel_4;
input 	Equal3;
input 	Equal31;
input 	Equal4;
output 	saved_grant_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	src4_valid;
input 	src4_valid1;
input 	last_channel_4;
input 	src4_valid2;
output 	src_valid;
output 	src_valid1;
output 	src_payload_0;
output 	src_data_78;
output 	src_data_79;
output 	src_data_35;
output 	src_data_34;
output 	src_data_33;
output 	src_data_32;
input 	Selector3;
input 	Selector10;
input 	Selector4;
input 	Selector11;
output 	src_payload;
output 	src_data_73;
output 	src_data_72;
output 	src_payload1;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
input 	nxt_in_ready2;
input 	src4_valid3;
output 	src_data_92;
output 	src_data_93;
output 	src_data_94;
output 	src_data_95;
output 	src_data_96;
output 	src_data_97;
output 	src_data_98;
output 	src_data_99;
output 	src_data_100;
output 	src_data_101;
output 	src_data_102;
output 	src_data_103;
output 	src_data_77;
input 	Selector5;
input 	Selector12;
output 	src_data_71;
input 	Selector6;
input 	nxt_out_burstwrap_0;
output 	src_data_70;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \arb|grant[0]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


terminal_qsys_altera_merlin_arbitrator_3 arb(
	.src_channel_4(src_channel_4),
	.Equal3(Equal3),
	.Equal31(Equal31),
	.Equal4(Equal4),
	.reset(altera_reset_synchronizer_int_chain_out),
	.src4_valid(src4_valid),
	.src4_valid1(src4_valid1),
	.src4_valid2(src4_valid2),
	.grant_1(\arb|grant[1]~0_combout ),
	.src_valid(src_valid),
	.src_valid1(src_valid1),
	.src_payload_0(src_payload_0),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_0(\arb|grant[0]~1_combout ),
	.nxt_in_ready(nxt_in_ready2),
	.src4_valid3(src4_valid3),
	.clk(clk_clk));

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cyclonev_lcell_comb \src_valid~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!saved_grant_1),
	.datac(!has_pending_responses),
	.datad(!src_channel_4),
	.datae(!last_channel_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~0 .extended_lut = "off";
defparam \src_valid~0 .lut_mask = 64'h0010001100100011;
defparam \src_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src_valid~1 (
	.dataa(!saved_grant_0),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(!Equal4),
	.datae(!src4_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_valid~1 .extended_lut = "off";
defparam \src_valid~1 .lut_mask = 64'h0000544400005444;
defparam \src_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload[0] (
	.dataa(!h2f_lw_WLAST_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h3737373737373737;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[78] (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!h2f_lw_AWSIZE_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_78),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[78] .extended_lut = "off";
defparam \src_data[78] .lut_mask = 64'h0537053705370537;
defparam \src_data[78] .shared_arith = "off";

cyclonev_lcell_comb \src_data[79] (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!h2f_lw_AWSIZE_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_79),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[79] .extended_lut = "off";
defparam \src_data[79] .lut_mask = 64'h0537053705370537;
defparam \src_data[79] .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!h2f_lw_WSTRB_3),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h3737373737373737;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!h2f_lw_WSTRB_2),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h3737373737373737;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!h2f_lw_WSTRB_1),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h3737373737373737;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!h2f_lw_WSTRB_0),
	.datab(!saved_grant_1),
	.datac(!saved_grant_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h3737373737373737;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_WDATA_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[73] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector3),
	.datad(!Selector10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_73),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[73] .extended_lut = "off";
defparam \src_data[73] .lut_mask = 64'h3075307530753075;
defparam \src_data[73] .shared_arith = "off";

cyclonev_lcell_comb \src_data[72] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector4),
	.datad(!Selector11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_72),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[72] .extended_lut = "off";
defparam \src_data[72] .lut_mask = 64'h3075307530753075;
defparam \src_data[72] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_WDATA_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_WDATA_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!h2f_lw_WDATA_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h1111111111111111;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!h2f_lw_WDATA_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h1111111111111111;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!h2f_lw_WDATA_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h1111111111111111;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!h2f_lw_WDATA_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h1111111111111111;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!h2f_lw_WDATA_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h1111111111111111;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!h2f_lw_WDATA_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h1111111111111111;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!h2f_lw_WDATA_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h1111111111111111;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!h2f_lw_ARID_0),
	.datab(!h2f_lw_AWID_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'h0537053705370537;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!h2f_lw_ARID_1),
	.datab(!h2f_lw_AWID_1),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'h0537053705370537;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!h2f_lw_ARID_2),
	.datab(!h2f_lw_AWID_2),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'h0537053705370537;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!h2f_lw_ARID_3),
	.datab(!h2f_lw_AWID_3),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'h0537053705370537;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!h2f_lw_ARID_4),
	.datab(!h2f_lw_AWID_4),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'h0537053705370537;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!h2f_lw_ARID_5),
	.datab(!h2f_lw_AWID_5),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'h0537053705370537;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!h2f_lw_ARID_6),
	.datab(!h2f_lw_AWID_6),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'h0537053705370537;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!h2f_lw_ARID_7),
	.datab(!h2f_lw_AWID_7),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'h0537053705370537;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[100] (
	.dataa(!h2f_lw_ARID_8),
	.datab(!h2f_lw_AWID_8),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_100),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100] .extended_lut = "off";
defparam \src_data[100] .lut_mask = 64'h0537053705370537;
defparam \src_data[100] .shared_arith = "off";

cyclonev_lcell_comb \src_data[101] (
	.dataa(!h2f_lw_ARID_9),
	.datab(!h2f_lw_AWID_9),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101] .extended_lut = "off";
defparam \src_data[101] .lut_mask = 64'h0537053705370537;
defparam \src_data[101] .shared_arith = "off";

cyclonev_lcell_comb \src_data[102] (
	.dataa(!h2f_lw_ARID_10),
	.datab(!h2f_lw_AWID_10),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102] .extended_lut = "off";
defparam \src_data[102] .lut_mask = 64'h0537053705370537;
defparam \src_data[102] .shared_arith = "off";

cyclonev_lcell_comb \src_data[103] (
	.dataa(!h2f_lw_ARID_11),
	.datab(!h2f_lw_AWID_11),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103] .extended_lut = "off";
defparam \src_data[103] .lut_mask = 64'h0537053705370537;
defparam \src_data[103] .shared_arith = "off";

cyclonev_lcell_comb \src_data[77] (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!h2f_lw_AWSIZE_0),
	.datac(!saved_grant_1),
	.datad(!saved_grant_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_77),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[77] .extended_lut = "off";
defparam \src_data[77] .lut_mask = 64'h0537053705370537;
defparam \src_data[77] .shared_arith = "off";

cyclonev_lcell_comb \src_data[71] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector5),
	.datad(!Selector12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_71),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[71] .extended_lut = "off";
defparam \src_data[71] .lut_mask = 64'h3075307530753075;
defparam \src_data[71] .shared_arith = "off";

cyclonev_lcell_comb \src_data[70] (
	.dataa(!saved_grant_1),
	.datab(!saved_grant_0),
	.datac(!Selector6),
	.datad(!nxt_out_burstwrap_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_70),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[70] .extended_lut = "off";
defparam \src_data[70] .lut_mask = 64'h3075307530753075;
defparam \src_data[70] .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!nxt_in_ready1),
	.datab(!nxt_in_ready),
	.datac(!src_valid),
	.datad(!src_valid1),
	.datae(!src_payload_0),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hF000F77700000777;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_merlin_arbitrator_3 (
	src_channel_4,
	Equal3,
	Equal31,
	Equal4,
	reset,
	src4_valid,
	src4_valid1,
	src4_valid2,
	grant_1,
	src_valid,
	src_valid1,
	src_payload_0,
	packet_in_progress,
	grant_0,
	nxt_in_ready,
	src4_valid3,
	clk)/* synthesis synthesis_greybox=0 */;
input 	src_channel_4;
input 	Equal3;
input 	Equal31;
input 	Equal4;
input 	reset;
input 	src4_valid;
input 	src4_valid1;
input 	src4_valid2;
output 	grant_1;
input 	src_valid;
input 	src_valid1;
input 	src_payload_0;
input 	packet_in_progress;
output 	grant_0;
input 	nxt_in_ready;
input 	src4_valid3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg[0]~2_combout ;
wire \top_priority_reg[0]~q ;


cyclonev_lcell_comb \grant[1]~0 (
	.dataa(!src4_valid),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!src4_valid1),
	.datae(!src4_valid2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~0 .extended_lut = "off";
defparam \grant[1]~0 .lut_mask = 64'h0000F3B30000F3B3;
defparam \grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[0]~1 (
	.dataa(!src4_valid),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!src4_valid1),
	.datae(!src4_valid2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~1 .extended_lut = "off";
defparam \grant[0]~1 .lut_mask = 64'h0051005000510050;
defparam \grant[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!src_channel_4),
	.datab(!Equal3),
	.datac(!Equal31),
	.datad(!Equal4),
	.datae(!src4_valid1),
	.dataf(!src4_valid3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'h0000FCCC5555FDDD;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!nxt_in_ready),
	.datab(!src_valid),
	.datac(!src_valid1),
	.datad(!src_payload_0),
	.datae(!packet_in_progress),
	.dataf(!\top_priority_reg[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'h00000000C0EA002A;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cyclonev_lcell_comb \top_priority_reg[0]~2 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~2 .extended_lut = "off";
defparam \top_priority_reg[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~2 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~1_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_cmd_mux_5 (
	h2f_lw_ARVALID_0,
	h2f_lw_ARSIZE_0,
	h2f_lw_ARSIZE_1,
	h2f_lw_ARSIZE_2,
	Equal5,
	saved_grant_1,
	nxt_in_ready,
	nxt_in_ready1,
	has_pending_responses,
	altera_reset_synchronizer_int_chain_out,
	last_channel_5,
	last_cycle,
	src_payload,
	src_payload1,
	src_payload2,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARVALID_0;
input 	h2f_lw_ARSIZE_0;
input 	h2f_lw_ARSIZE_1;
input 	h2f_lw_ARSIZE_2;
input 	Equal5;
output 	saved_grant_1;
input 	nxt_in_ready;
input 	nxt_in_ready1;
input 	has_pending_responses;
input 	altera_reset_synchronizer_int_chain_out;
input 	last_channel_5;
output 	last_cycle;
output 	src_payload;
output 	src_payload1;
output 	src_payload2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \saved_grant[1]~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \saved_grant[1]~1_combout ;


dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\saved_grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \last_cycle~0 (
	.dataa(!saved_grant_1),
	.datab(!\saved_grant[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(last_cycle),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_cycle~0 .extended_lut = "off";
defparam \last_cycle~0 .lut_mask = 64'h1111111111111111;
defparam \last_cycle~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!h2f_lw_ARSIZE_0),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h1111111111111111;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!h2f_lw_ARSIZE_2),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h1111111111111111;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!h2f_lw_ARSIZE_1),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h1111111111111111;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \saved_grant[1]~0 (
	.dataa(!h2f_lw_ARVALID_0),
	.datab(!has_pending_responses),
	.datac(!last_channel_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~0 .extended_lut = "off";
defparam \saved_grant[1]~0 .lut_mask = 64'h4545454545454545;
defparam \saved_grant[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\saved_grant[1]~0_combout ),
	.datab(!saved_grant_1),
	.datac(!nxt_in_ready1),
	.datad(!nxt_in_ready),
	.datae(!\packet_in_progress~q ),
	.dataf(!Equal5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h0000FFFF0100EFEE;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \saved_grant[1]~1 (
	.dataa(!Equal5),
	.datab(!saved_grant_1),
	.datac(gnd),
	.datad(!\saved_grant[1]~0_combout ),
	.datae(!\packet_in_progress~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\saved_grant[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \saved_grant[1]~1 .extended_lut = "off";
defparam \saved_grant[1]~1 .lut_mask = 64'h0055333300553333;
defparam \saved_grant[1]~1 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_router (
	h2f_lw_AWADDR_4,
	h2f_lw_AWADDR_5,
	h2f_lw_AWADDR_6,
	h2f_lw_AWADDR_7,
	h2f_lw_AWADDR_8,
	h2f_lw_AWADDR_9,
	h2f_lw_AWADDR_10,
	h2f_lw_AWADDR_11,
	h2f_lw_AWADDR_12,
	h2f_lw_AWADDR_13,
	h2f_lw_AWADDR_14,
	h2f_lw_AWADDR_15,
	address_burst_7,
	address_burst_6,
	address_burst_9,
	address_burst_8,
	address_burst_11,
	address_burst_10,
	address_burst_15,
	address_burst_14,
	address_burst_13,
	address_burst_12,
	sop_enable,
	address_burst_5,
	address_burst_4,
	Equal3,
	out_data_18,
	out_data_17,
	out_data_16,
	Equal31,
	Equal4,
	Equal32,
	Equal41)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_AWADDR_4;
input 	h2f_lw_AWADDR_5;
input 	h2f_lw_AWADDR_6;
input 	h2f_lw_AWADDR_7;
input 	h2f_lw_AWADDR_8;
input 	h2f_lw_AWADDR_9;
input 	h2f_lw_AWADDR_10;
input 	h2f_lw_AWADDR_11;
input 	h2f_lw_AWADDR_12;
input 	h2f_lw_AWADDR_13;
input 	h2f_lw_AWADDR_14;
input 	h2f_lw_AWADDR_15;
input 	address_burst_7;
input 	address_burst_6;
input 	address_burst_9;
input 	address_burst_8;
input 	address_burst_11;
input 	address_burst_10;
input 	address_burst_15;
input 	address_burst_14;
input 	address_burst_13;
input 	address_burst_12;
input 	sop_enable;
input 	address_burst_5;
input 	address_burst_4;
output 	Equal3;
input 	out_data_18;
input 	out_data_17;
input 	out_data_16;
output 	Equal31;
output 	Equal4;
output 	Equal32;
output 	Equal41;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal3~0_combout ;
wire \Equal3~1_combout ;
wire \Equal3~2_combout ;
wire \Equal3~3_combout ;
wire \Equal3~4_combout ;
wire \Equal3~5_combout ;


cyclonev_lcell_comb \Equal3~6 (
	.dataa(!\Equal3~0_combout ),
	.datab(!\Equal3~1_combout ),
	.datac(!\Equal3~2_combout ),
	.datad(!\Equal3~3_combout ),
	.datae(!\Equal3~4_combout ),
	.dataf(!\Equal3~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~6 .extended_lut = "off";
defparam \Equal3~6 .lut_mask = 64'h0000000000000001;
defparam \Equal3~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~7 (
	.dataa(!out_data_18),
	.datab(!out_data_17),
	.datac(!out_data_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~7 .extended_lut = "off";
defparam \Equal3~7 .lut_mask = 64'h0202020202020202;
defparam \Equal3~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!out_data_18),
	.datab(!out_data_17),
	.datac(!out_data_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h4040404040404040;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~8 (
	.dataa(!Equal3),
	.datab(!Equal31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~8 .extended_lut = "off";
defparam \Equal3~8 .lut_mask = 64'h1111111111111111;
defparam \Equal3~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!Equal3),
	.datab(!Equal4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal41),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h1111111111111111;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!h2f_lw_AWADDR_4),
	.datab(!h2f_lw_AWADDR_5),
	.datac(!sop_enable),
	.datad(!address_burst_5),
	.datae(!address_burst_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h8F8080808F808080;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~1 (
	.dataa(!h2f_lw_AWADDR_6),
	.datab(!h2f_lw_AWADDR_7),
	.datac(!sop_enable),
	.datad(!address_burst_7),
	.datae(!address_burst_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~1 .extended_lut = "off";
defparam \Equal3~1 .lut_mask = 64'h8F8080808F808080;
defparam \Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~2 (
	.dataa(!h2f_lw_AWADDR_8),
	.datab(!h2f_lw_AWADDR_9),
	.datac(!sop_enable),
	.datad(!address_burst_9),
	.datae(!address_burst_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~2 .extended_lut = "off";
defparam \Equal3~2 .lut_mask = 64'h8F8080808F808080;
defparam \Equal3~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~3 (
	.dataa(!h2f_lw_AWADDR_10),
	.datab(!h2f_lw_AWADDR_11),
	.datac(!sop_enable),
	.datad(!address_burst_11),
	.datae(!address_burst_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~3 .extended_lut = "off";
defparam \Equal3~3 .lut_mask = 64'h8F8080808F808080;
defparam \Equal3~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~4 (
	.dataa(!h2f_lw_AWADDR_14),
	.datab(!h2f_lw_AWADDR_15),
	.datac(!sop_enable),
	.datad(!address_burst_15),
	.datae(!address_burst_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~4 .extended_lut = "off";
defparam \Equal3~4 .lut_mask = 64'h8F8080808F808080;
defparam \Equal3~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~5 (
	.dataa(!h2f_lw_AWADDR_12),
	.datab(!h2f_lw_AWADDR_13),
	.datac(!sop_enable),
	.datad(!address_burst_13),
	.datae(!address_burst_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~5 .extended_lut = "off";
defparam \Equal3~5 .lut_mask = 64'h8F8080808F808080;
defparam \Equal3~5 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_router_1 (
	h2f_lw_ARADDR_3,
	h2f_lw_ARADDR_4,
	h2f_lw_ARADDR_5,
	h2f_lw_ARADDR_6,
	h2f_lw_ARADDR_7,
	h2f_lw_ARADDR_8,
	h2f_lw_ARADDR_9,
	h2f_lw_ARADDR_10,
	h2f_lw_ARADDR_11,
	h2f_lw_ARADDR_12,
	h2f_lw_ARADDR_13,
	h2f_lw_ARADDR_14,
	h2f_lw_ARADDR_15,
	h2f_lw_ARADDR_16,
	h2f_lw_ARADDR_17,
	h2f_lw_ARADDR_18,
	Equal1,
	Equal11,
	Equal5,
	src_channel_4,
	Equal4,
	Equal41,
	Equal12,
	Equal3,
	src_channel_41,
	src_data_90,
	src_data_91,
	Equal13,
	Equal2)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_ARADDR_3;
input 	h2f_lw_ARADDR_4;
input 	h2f_lw_ARADDR_5;
input 	h2f_lw_ARADDR_6;
input 	h2f_lw_ARADDR_7;
input 	h2f_lw_ARADDR_8;
input 	h2f_lw_ARADDR_9;
input 	h2f_lw_ARADDR_10;
input 	h2f_lw_ARADDR_11;
input 	h2f_lw_ARADDR_12;
input 	h2f_lw_ARADDR_13;
input 	h2f_lw_ARADDR_14;
input 	h2f_lw_ARADDR_15;
input 	h2f_lw_ARADDR_16;
input 	h2f_lw_ARADDR_17;
input 	h2f_lw_ARADDR_18;
output 	Equal1;
output 	Equal11;
output 	Equal5;
output 	src_channel_4;
output 	Equal4;
output 	Equal41;
output 	Equal12;
output 	Equal3;
output 	src_channel_41;
output 	src_data_90;
output 	src_data_91;
output 	Equal13;
output 	Equal2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!h2f_lw_ARADDR_4),
	.datab(!h2f_lw_ARADDR_5),
	.datac(!h2f_lw_ARADDR_6),
	.datad(!h2f_lw_ARADDR_7),
	.datae(!h2f_lw_ARADDR_8),
	.dataf(!h2f_lw_ARADDR_9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h8000000000000000;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!h2f_lw_ARADDR_10),
	.datab(!h2f_lw_ARADDR_11),
	.datac(!h2f_lw_ARADDR_12),
	.datad(!h2f_lw_ARADDR_13),
	.datae(!h2f_lw_ARADDR_14),
	.dataf(!h2f_lw_ARADDR_15),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'h8000000000000000;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!h2f_lw_ARADDR_18),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'h0000000200000002;
defparam \Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[4]~0 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!h2f_lw_ARADDR_16),
	.datac(!h2f_lw_ARADDR_17),
	.datad(!h2f_lw_ARADDR_18),
	.datae(!Equal1),
	.dataf(!Equal11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[4]~0 .extended_lut = "off";
defparam \src_channel[4]~0 .lut_mask = 64'h000000000000230C;
defparam \src_channel[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!h2f_lw_ARADDR_17),
	.datab(!h2f_lw_ARADDR_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h2222222222222222;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!Equal4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal41),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h0002000200020002;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~2 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~2 .extended_lut = "off";
defparam \Equal1~2 .lut_mask = 64'h4444444444444444;
defparam \Equal1~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!h2f_lw_ARADDR_17),
	.datab(!Equal1),
	.datac(!Equal11),
	.datad(!Equal12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h0001000100010001;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \src_channel[4]~1 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!h2f_lw_ARADDR_16),
	.datac(!h2f_lw_ARADDR_17),
	.datad(!h2f_lw_ARADDR_18),
	.datae(!Equal1),
	.dataf(!Equal11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_channel_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_channel[4]~1 .extended_lut = "off";
defparam \src_channel[4]~1 .lut_mask = 64'hFFFFFFFFFFFFD033;
defparam \src_channel[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[90]~0 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!h2f_lw_ARADDR_18),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_90),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[90]~0 .extended_lut = "off";
defparam \src_data[90]~0 .lut_mask = 64'hFFFFFFC5FFFFFFC5;
defparam \src_data[90]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[91]~1 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(gnd),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_91),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[91]~1 .extended_lut = "off";
defparam \src_data[91]~1 .lut_mask = 64'h0000002200000022;
defparam \src_data[91]~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~3 (
	.dataa(!h2f_lw_ARADDR_3),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!Equal1),
	.datad(!Equal11),
	.datae(!Equal12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~3 .extended_lut = "off";
defparam \Equal1~3 .lut_mask = 64'h0000000800000008;
defparam \Equal1~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!h2f_lw_ARADDR_16),
	.datab(!h2f_lw_ARADDR_17),
	.datac(!h2f_lw_ARADDR_18),
	.datad(!Equal1),
	.datae(!Equal11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h0000002000000020;
defparam \Equal2~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_demux_2 (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_59_0),
	.datad(!mem_57_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_demux_3 (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_59_0),
	.datad(!mem_57_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_demux_4 (
	h2f_lw_BREADY_0,
	h2f_lw_RREADY_0,
	read_latency_shift_reg_0,
	mem_used_0,
	mem_116_0,
	mem_used_01,
	mem_59_0,
	mem_57_0,
	src0_valid1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=0 */;
input 	h2f_lw_BREADY_0;
input 	h2f_lw_RREADY_0;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	mem_116_0;
input 	mem_used_01;
input 	mem_59_0;
input 	mem_57_0;
output 	src0_valid1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb src0_valid(
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam src0_valid.extended_lut = "off";
defparam src0_valid.lut_mask = 64'h0000777F00000000;
defparam src0_valid.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_116_0),
	.datad(!mem_used_01),
	.datae(!mem_59_0),
	.dataf(!mem_57_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h8880FFFF88808880;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!h2f_lw_BREADY_0),
	.datab(!h2f_lw_RREADY_0),
	.datac(!mem_59_0),
	.datad(!mem_57_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h3533353335333533;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_mux (
	src0_valid,
	src0_valid1,
	src0_valid2,
	WideOr11,
	mem_92_0,
	mem_92_01,
	mem_92_02,
	src_payload,
	mem_93_0,
	mem_93_01,
	mem_93_02,
	src_payload1,
	mem_94_0,
	mem_94_01,
	mem_94_02,
	src_payload2,
	mem_95_0,
	mem_95_01,
	mem_95_02,
	src_payload3,
	mem_96_0,
	mem_96_01,
	mem_96_02,
	src_payload4,
	mem_97_0,
	mem_97_01,
	mem_97_02,
	src_payload5,
	mem_98_0,
	mem_98_01,
	mem_98_02,
	src_payload6,
	mem_99_0,
	mem_99_01,
	mem_99_02,
	src_payload7,
	mem_100_0,
	mem_100_01,
	mem_100_02,
	src_payload8,
	mem_101_0,
	mem_101_01,
	mem_101_02,
	src_payload9,
	mem_102_0,
	mem_102_01,
	mem_102_02,
	src_payload10,
	mem_103_0,
	mem_103_01,
	mem_103_02,
	src_payload11)/* synthesis synthesis_greybox=0 */;
input 	src0_valid;
input 	src0_valid1;
input 	src0_valid2;
output 	WideOr11;
input 	mem_92_0;
input 	mem_92_01;
input 	mem_92_02;
output 	src_payload;
input 	mem_93_0;
input 	mem_93_01;
input 	mem_93_02;
output 	src_payload1;
input 	mem_94_0;
input 	mem_94_01;
input 	mem_94_02;
output 	src_payload2;
input 	mem_95_0;
input 	mem_95_01;
input 	mem_95_02;
output 	src_payload3;
input 	mem_96_0;
input 	mem_96_01;
input 	mem_96_02;
output 	src_payload4;
input 	mem_97_0;
input 	mem_97_01;
input 	mem_97_02;
output 	src_payload5;
input 	mem_98_0;
input 	mem_98_01;
input 	mem_98_02;
output 	src_payload6;
input 	mem_99_0;
input 	mem_99_01;
input 	mem_99_02;
output 	src_payload7;
input 	mem_100_0;
input 	mem_100_01;
input 	mem_100_02;
output 	src_payload8;
input 	mem_101_0;
input 	mem_101_01;
input 	mem_101_02;
output 	src_payload9;
input 	mem_102_0;
input 	mem_102_01;
input 	mem_102_02;
output 	src_payload10;
input 	mem_103_0;
input 	mem_103_01;
input 	mem_103_02;
output 	src_payload11;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb WideOr1(
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_92_0),
	.datae(!mem_92_01),
	.dataf(!mem_92_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_93_0),
	.datae(!mem_93_01),
	.dataf(!mem_93_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_94_0),
	.datae(!mem_94_01),
	.dataf(!mem_94_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_95_0),
	.datae(!mem_95_01),
	.dataf(!mem_95_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_96_0),
	.datae(!mem_96_01),
	.dataf(!mem_96_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_97_0),
	.datae(!mem_97_01),
	.dataf(!mem_97_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_98_0),
	.datae(!mem_98_01),
	.dataf(!mem_98_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_99_0),
	.datae(!mem_99_01),
	.dataf(!mem_99_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_100_0),
	.datae(!mem_100_01),
	.dataf(!mem_100_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_101_0),
	.datae(!mem_101_01),
	.dataf(!mem_101_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_102_0),
	.datae(!mem_102_01),
	.dataf(!mem_102_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!src0_valid2),
	.datad(!mem_103_0),
	.datae(!mem_103_01),
	.dataf(!mem_103_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h005533770F5F3F7F;
defparam \src_payload~11 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_mm_interconnect_0_rsp_mux_1 (
	in_ready_hold,
	mem_57_0,
	mem_57_01,
	mem_57_02,
	comb,
	src1_valid,
	mem_117_0,
	last_packet_beat,
	last_packet_beat1,
	comb1,
	src1_valid1,
	mem_117_01,
	last_packet_beat2,
	last_packet_beat3,
	comb2,
	src1_valid2,
	mem_117_02,
	last_packet_beat4,
	last_packet_beat5,
	mem_117_03,
	read_latency_shift_reg_0,
	mem_used_0,
	empty,
	mem_57_03,
	mem_used_01,
	last_packet_beat6,
	last_packet_beat7,
	mem_117_04,
	read_latency_shift_reg_01,
	mem_used_02,
	empty1,
	mem_57_04,
	mem_used_03,
	last_packet_beat8,
	last_packet_beat9,
	mem_117_05,
	read_latency_shift_reg_02,
	mem_used_04,
	empty2,
	mem_57_05,
	mem_used_05,
	last_packet_beat10,
	last_packet_beat11,
	src_payload_0,
	WideOr11,
	mem_92_0,
	mem_92_01,
	mem_92_02,
	mem_93_0,
	mem_93_01,
	mem_93_02,
	mem_94_0,
	mem_94_01,
	mem_94_02,
	mem_95_0,
	mem_95_01,
	mem_95_02,
	mem_96_0,
	mem_96_01,
	mem_96_02,
	mem_97_0,
	mem_97_01,
	mem_97_02,
	mem_98_0,
	mem_98_01,
	mem_98_02,
	mem_99_0,
	mem_99_01,
	mem_99_02,
	mem_100_0,
	mem_100_01,
	mem_100_02,
	mem_101_0,
	mem_101_01,
	mem_101_02,
	mem_102_0,
	mem_102_01,
	mem_102_02,
	mem_103_0,
	mem_103_01,
	mem_103_02,
	av_readdata_pre_0,
	always4,
	mem_0_0,
	av_readdata_pre_01,
	always41,
	mem_0_01,
	av_readdata_pre_02,
	always42,
	mem_0_02,
	mem_0_03,
	av_readdata_pre_03,
	mem_0_04,
	av_readdata_pre_04,
	src_data_0,
	av_readdata_pre_1,
	mem_1_0,
	av_readdata_pre_11,
	mem_1_01,
	av_readdata_pre_12,
	mem_1_02,
	mem_1_03,
	av_readdata_pre_13,
	mem_1_04,
	av_readdata_pre_14,
	src_data_1,
	av_readdata_pre_2,
	mem_2_0,
	av_readdata_pre_21,
	mem_2_01,
	av_readdata_pre_22,
	mem_2_02,
	mem_2_03,
	av_readdata_pre_23,
	mem_11_0,
	av_readdata_pre_30,
	mem_2_04,
	av_readdata_pre_24,
	src_data_2,
	av_readdata_pre_3,
	mem_3_0,
	av_readdata_pre_31,
	mem_3_01,
	av_readdata_pre_32,
	mem_3_02,
	mem_3_03,
	av_readdata_pre_33,
	mem_3_04,
	av_readdata_pre_34,
	src_data_3,
	av_readdata_pre_4,
	mem_4_0,
	av_readdata_pre_41,
	mem_4_01,
	av_readdata_pre_42,
	mem_4_02,
	mem_4_03,
	av_readdata_pre_43,
	mem_4_04,
	av_readdata_pre_44,
	src_data_4,
	av_readdata_pre_5,
	mem_5_0,
	av_readdata_pre_51,
	mem_5_01,
	av_readdata_pre_52,
	mem_5_02,
	mem_5_03,
	av_readdata_pre_53,
	mem_5_04,
	av_readdata_pre_54,
	src_data_5,
	av_readdata_pre_6,
	mem_6_0,
	av_readdata_pre_61,
	mem_6_01,
	av_readdata_pre_62,
	mem_6_02,
	mem_6_03,
	av_readdata_pre_63,
	mem_6_04,
	av_readdata_pre_64,
	src_data_6,
	av_readdata_pre_7,
	mem_7_0,
	av_readdata_pre_71,
	mem_7_01,
	av_readdata_pre_72,
	mem_7_02,
	mem_7_03,
	av_readdata_pre_73,
	mem_10_0,
	mem_7_04,
	av_readdata_pre_74,
	src_data_7,
	av_readdata_pre_8,
	mem_8_0,
	av_readdata_pre_81,
	mem_8_01,
	av_readdata_pre_82,
	mem_8_02,
	mem_8_03,
	av_readdata_pre_83,
	mem_8_04,
	av_readdata_pre_84,
	src_data_8,
	av_readdata_pre_9,
	av_readdata_pre_91,
	mem_9_0,
	av_readdata_pre_92,
	mem_9_01,
	av_readdata_pre_93,
	mem_9_02,
	mem_9_03,
	av_readdata_pre_94,
	mem_9_04,
	src_data_9,
	av_readdata_pre_10,
	mem_10_01,
	av_readdata_pre_101,
	mem_10_02,
	mem_10_03,
	av_readdata_pre_102,
	src_payload,
	av_readdata_pre_111,
	mem_11_01,
	av_readdata_pre_112,
	mem_11_02,
	mem_11_03,
	av_readdata_pre_113,
	src_payload1,
	av_readdata_pre_121,
	mem_12_0,
	av_readdata_pre_122,
	mem_12_01,
	mem_12_02,
	av_readdata_pre_123,
	src_payload2,
	av_readdata_pre_131,
	mem_13_0,
	av_readdata_pre_132,
	mem_13_01,
	mem_13_02,
	av_readdata_pre_133,
	src_payload3,
	av_readdata_pre_141,
	mem_14_0,
	av_readdata_pre_142,
	mem_14_01,
	mem_14_02,
	av_readdata_pre_143,
	src_payload4,
	av_readdata_pre_15,
	mem_15_0,
	av_readdata_pre_151,
	mem_15_01,
	mem_15_02,
	av_readdata_pre_152,
	src_payload5,
	av_readdata_pre_16,
	mem_16_0,
	av_readdata_pre_161,
	mem_16_01,
	mem_16_02,
	av_readdata_pre_162,
	src_payload6,
	av_readdata_pre_17,
	mem_17_0,
	av_readdata_pre_171,
	mem_17_01,
	mem_17_02,
	av_readdata_pre_172,
	src_payload7,
	av_readdata_pre_18,
	mem_18_0,
	av_readdata_pre_181,
	mem_18_01,
	mem_18_02,
	av_readdata_pre_182,
	src_payload8,
	av_readdata_pre_19,
	mem_19_0,
	av_readdata_pre_191,
	mem_19_01,
	mem_19_02,
	av_readdata_pre_192,
	src_payload9,
	av_readdata_pre_20,
	mem_20_0,
	av_readdata_pre_201,
	mem_20_01,
	mem_20_02,
	av_readdata_pre_202,
	src_payload10,
	av_readdata_pre_211,
	mem_21_0,
	av_readdata_pre_212,
	mem_21_01,
	mem_21_02,
	av_readdata_pre_213,
	src_payload11,
	av_readdata_pre_221,
	mem_22_0,
	av_readdata_pre_222,
	mem_22_01,
	mem_22_02,
	av_readdata_pre_223,
	src_payload12,
	av_readdata_pre_231,
	mem_23_0,
	av_readdata_pre_232,
	mem_23_01,
	mem_23_02,
	av_readdata_pre_233,
	src_payload13,
	av_readdata_pre_241,
	mem_24_0,
	av_readdata_pre_242,
	mem_24_01,
	mem_24_02,
	av_readdata_pre_243,
	src_payload14,
	av_readdata_pre_25,
	mem_25_0,
	av_readdata_pre_251,
	mem_25_01,
	mem_25_02,
	av_readdata_pre_252,
	src_payload15,
	av_readdata_pre_26,
	mem_26_0,
	av_readdata_pre_261,
	mem_26_01,
	mem_26_02,
	av_readdata_pre_262,
	src_payload16,
	av_readdata_pre_27,
	mem_27_0,
	av_readdata_pre_271,
	mem_27_01,
	mem_27_02,
	av_readdata_pre_272,
	src_payload17,
	av_readdata_pre_28,
	mem_28_0,
	av_readdata_pre_281,
	mem_28_01,
	mem_28_02,
	av_readdata_pre_282,
	src_payload18,
	av_readdata_pre_29,
	mem_29_0,
	av_readdata_pre_291,
	mem_29_01,
	mem_29_02,
	av_readdata_pre_292,
	src_payload19,
	av_readdata_pre_301,
	mem_30_0,
	av_readdata_pre_302,
	mem_30_01,
	mem_30_02,
	av_readdata_pre_303,
	src_payload20,
	av_readdata_pre_311,
	mem_31_0,
	av_readdata_pre_312,
	mem_31_01,
	mem_31_02,
	av_readdata_pre_313,
	src_payload21,
	mem_92_03,
	mem_92_04,
	mem_92_05,
	src_data_92,
	mem_93_03,
	mem_93_04,
	mem_93_05,
	src_data_93,
	mem_94_03,
	mem_94_04,
	mem_94_05,
	src_data_94,
	mem_95_03,
	mem_95_04,
	mem_95_05,
	src_data_95,
	mem_96_03,
	mem_96_04,
	mem_96_05,
	src_data_96,
	mem_97_03,
	mem_97_04,
	mem_97_05,
	src_data_97,
	mem_98_03,
	mem_98_04,
	mem_98_05,
	src_data_98,
	mem_99_03,
	mem_99_04,
	mem_99_05,
	src_data_99,
	mem_100_03,
	mem_100_04,
	mem_100_05,
	src_data_100,
	mem_101_03,
	mem_101_04,
	mem_101_05,
	src_data_101,
	mem_102_03,
	mem_102_04,
	mem_102_05,
	src_data_102,
	mem_103_03,
	mem_103_04,
	mem_103_05,
	src_data_103,
	src_payload22)/* synthesis synthesis_greybox=0 */;
input 	in_ready_hold;
input 	mem_57_0;
input 	mem_57_01;
input 	mem_57_02;
input 	comb;
input 	src1_valid;
input 	mem_117_0;
input 	last_packet_beat;
input 	last_packet_beat1;
input 	comb1;
input 	src1_valid1;
input 	mem_117_01;
input 	last_packet_beat2;
input 	last_packet_beat3;
input 	comb2;
input 	src1_valid2;
input 	mem_117_02;
input 	last_packet_beat4;
input 	last_packet_beat5;
input 	mem_117_03;
input 	read_latency_shift_reg_0;
input 	mem_used_0;
input 	empty;
input 	mem_57_03;
input 	mem_used_01;
input 	last_packet_beat6;
input 	last_packet_beat7;
input 	mem_117_04;
input 	read_latency_shift_reg_01;
input 	mem_used_02;
input 	empty1;
input 	mem_57_04;
input 	mem_used_03;
input 	last_packet_beat8;
input 	last_packet_beat9;
input 	mem_117_05;
input 	read_latency_shift_reg_02;
input 	mem_used_04;
input 	empty2;
input 	mem_57_05;
input 	mem_used_05;
input 	last_packet_beat10;
input 	last_packet_beat11;
output 	src_payload_0;
output 	WideOr11;
input 	mem_92_0;
input 	mem_92_01;
input 	mem_92_02;
input 	mem_93_0;
input 	mem_93_01;
input 	mem_93_02;
input 	mem_94_0;
input 	mem_94_01;
input 	mem_94_02;
input 	mem_95_0;
input 	mem_95_01;
input 	mem_95_02;
input 	mem_96_0;
input 	mem_96_01;
input 	mem_96_02;
input 	mem_97_0;
input 	mem_97_01;
input 	mem_97_02;
input 	mem_98_0;
input 	mem_98_01;
input 	mem_98_02;
input 	mem_99_0;
input 	mem_99_01;
input 	mem_99_02;
input 	mem_100_0;
input 	mem_100_01;
input 	mem_100_02;
input 	mem_101_0;
input 	mem_101_01;
input 	mem_101_02;
input 	mem_102_0;
input 	mem_102_01;
input 	mem_102_02;
input 	mem_103_0;
input 	mem_103_01;
input 	mem_103_02;
input 	av_readdata_pre_0;
input 	always4;
input 	mem_0_0;
input 	av_readdata_pre_01;
input 	always41;
input 	mem_0_01;
input 	av_readdata_pre_02;
input 	always42;
input 	mem_0_02;
input 	mem_0_03;
input 	av_readdata_pre_03;
input 	mem_0_04;
input 	av_readdata_pre_04;
output 	src_data_0;
input 	av_readdata_pre_1;
input 	mem_1_0;
input 	av_readdata_pre_11;
input 	mem_1_01;
input 	av_readdata_pre_12;
input 	mem_1_02;
input 	mem_1_03;
input 	av_readdata_pre_13;
input 	mem_1_04;
input 	av_readdata_pre_14;
output 	src_data_1;
input 	av_readdata_pre_2;
input 	mem_2_0;
input 	av_readdata_pre_21;
input 	mem_2_01;
input 	av_readdata_pre_22;
input 	mem_2_02;
input 	mem_2_03;
input 	av_readdata_pre_23;
input 	mem_11_0;
input 	av_readdata_pre_30;
input 	mem_2_04;
input 	av_readdata_pre_24;
output 	src_data_2;
input 	av_readdata_pre_3;
input 	mem_3_0;
input 	av_readdata_pre_31;
input 	mem_3_01;
input 	av_readdata_pre_32;
input 	mem_3_02;
input 	mem_3_03;
input 	av_readdata_pre_33;
input 	mem_3_04;
input 	av_readdata_pre_34;
output 	src_data_3;
input 	av_readdata_pre_4;
input 	mem_4_0;
input 	av_readdata_pre_41;
input 	mem_4_01;
input 	av_readdata_pre_42;
input 	mem_4_02;
input 	mem_4_03;
input 	av_readdata_pre_43;
input 	mem_4_04;
input 	av_readdata_pre_44;
output 	src_data_4;
input 	av_readdata_pre_5;
input 	mem_5_0;
input 	av_readdata_pre_51;
input 	mem_5_01;
input 	av_readdata_pre_52;
input 	mem_5_02;
input 	mem_5_03;
input 	av_readdata_pre_53;
input 	mem_5_04;
input 	av_readdata_pre_54;
output 	src_data_5;
input 	av_readdata_pre_6;
input 	mem_6_0;
input 	av_readdata_pre_61;
input 	mem_6_01;
input 	av_readdata_pre_62;
input 	mem_6_02;
input 	mem_6_03;
input 	av_readdata_pre_63;
input 	mem_6_04;
input 	av_readdata_pre_64;
output 	src_data_6;
input 	av_readdata_pre_7;
input 	mem_7_0;
input 	av_readdata_pre_71;
input 	mem_7_01;
input 	av_readdata_pre_72;
input 	mem_7_02;
input 	mem_7_03;
input 	av_readdata_pre_73;
input 	mem_10_0;
input 	mem_7_04;
input 	av_readdata_pre_74;
output 	src_data_7;
input 	av_readdata_pre_8;
input 	mem_8_0;
input 	av_readdata_pre_81;
input 	mem_8_01;
input 	av_readdata_pre_82;
input 	mem_8_02;
input 	mem_8_03;
input 	av_readdata_pre_83;
input 	mem_8_04;
input 	av_readdata_pre_84;
output 	src_data_8;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
input 	mem_9_0;
input 	av_readdata_pre_92;
input 	mem_9_01;
input 	av_readdata_pre_93;
input 	mem_9_02;
input 	mem_9_03;
input 	av_readdata_pre_94;
input 	mem_9_04;
output 	src_data_9;
input 	av_readdata_pre_10;
input 	mem_10_01;
input 	av_readdata_pre_101;
input 	mem_10_02;
input 	mem_10_03;
input 	av_readdata_pre_102;
output 	src_payload;
input 	av_readdata_pre_111;
input 	mem_11_01;
input 	av_readdata_pre_112;
input 	mem_11_02;
input 	mem_11_03;
input 	av_readdata_pre_113;
output 	src_payload1;
input 	av_readdata_pre_121;
input 	mem_12_0;
input 	av_readdata_pre_122;
input 	mem_12_01;
input 	mem_12_02;
input 	av_readdata_pre_123;
output 	src_payload2;
input 	av_readdata_pre_131;
input 	mem_13_0;
input 	av_readdata_pre_132;
input 	mem_13_01;
input 	mem_13_02;
input 	av_readdata_pre_133;
output 	src_payload3;
input 	av_readdata_pre_141;
input 	mem_14_0;
input 	av_readdata_pre_142;
input 	mem_14_01;
input 	mem_14_02;
input 	av_readdata_pre_143;
output 	src_payload4;
input 	av_readdata_pre_15;
input 	mem_15_0;
input 	av_readdata_pre_151;
input 	mem_15_01;
input 	mem_15_02;
input 	av_readdata_pre_152;
output 	src_payload5;
input 	av_readdata_pre_16;
input 	mem_16_0;
input 	av_readdata_pre_161;
input 	mem_16_01;
input 	mem_16_02;
input 	av_readdata_pre_162;
output 	src_payload6;
input 	av_readdata_pre_17;
input 	mem_17_0;
input 	av_readdata_pre_171;
input 	mem_17_01;
input 	mem_17_02;
input 	av_readdata_pre_172;
output 	src_payload7;
input 	av_readdata_pre_18;
input 	mem_18_0;
input 	av_readdata_pre_181;
input 	mem_18_01;
input 	mem_18_02;
input 	av_readdata_pre_182;
output 	src_payload8;
input 	av_readdata_pre_19;
input 	mem_19_0;
input 	av_readdata_pre_191;
input 	mem_19_01;
input 	mem_19_02;
input 	av_readdata_pre_192;
output 	src_payload9;
input 	av_readdata_pre_20;
input 	mem_20_0;
input 	av_readdata_pre_201;
input 	mem_20_01;
input 	mem_20_02;
input 	av_readdata_pre_202;
output 	src_payload10;
input 	av_readdata_pre_211;
input 	mem_21_0;
input 	av_readdata_pre_212;
input 	mem_21_01;
input 	mem_21_02;
input 	av_readdata_pre_213;
output 	src_payload11;
input 	av_readdata_pre_221;
input 	mem_22_0;
input 	av_readdata_pre_222;
input 	mem_22_01;
input 	mem_22_02;
input 	av_readdata_pre_223;
output 	src_payload12;
input 	av_readdata_pre_231;
input 	mem_23_0;
input 	av_readdata_pre_232;
input 	mem_23_01;
input 	mem_23_02;
input 	av_readdata_pre_233;
output 	src_payload13;
input 	av_readdata_pre_241;
input 	mem_24_0;
input 	av_readdata_pre_242;
input 	mem_24_01;
input 	mem_24_02;
input 	av_readdata_pre_243;
output 	src_payload14;
input 	av_readdata_pre_25;
input 	mem_25_0;
input 	av_readdata_pre_251;
input 	mem_25_01;
input 	mem_25_02;
input 	av_readdata_pre_252;
output 	src_payload15;
input 	av_readdata_pre_26;
input 	mem_26_0;
input 	av_readdata_pre_261;
input 	mem_26_01;
input 	mem_26_02;
input 	av_readdata_pre_262;
output 	src_payload16;
input 	av_readdata_pre_27;
input 	mem_27_0;
input 	av_readdata_pre_271;
input 	mem_27_01;
input 	mem_27_02;
input 	av_readdata_pre_272;
output 	src_payload17;
input 	av_readdata_pre_28;
input 	mem_28_0;
input 	av_readdata_pre_281;
input 	mem_28_01;
input 	mem_28_02;
input 	av_readdata_pre_282;
output 	src_payload18;
input 	av_readdata_pre_29;
input 	mem_29_0;
input 	av_readdata_pre_291;
input 	mem_29_01;
input 	mem_29_02;
input 	av_readdata_pre_292;
output 	src_payload19;
input 	av_readdata_pre_301;
input 	mem_30_0;
input 	av_readdata_pre_302;
input 	mem_30_01;
input 	mem_30_02;
input 	av_readdata_pre_303;
output 	src_payload20;
input 	av_readdata_pre_311;
input 	mem_31_0;
input 	av_readdata_pre_312;
input 	mem_31_01;
input 	mem_31_02;
input 	av_readdata_pre_313;
output 	src_payload21;
input 	mem_92_03;
input 	mem_92_04;
input 	mem_92_05;
output 	src_data_92;
input 	mem_93_03;
input 	mem_93_04;
input 	mem_93_05;
output 	src_data_93;
input 	mem_94_03;
input 	mem_94_04;
input 	mem_94_05;
output 	src_data_94;
input 	mem_95_03;
input 	mem_95_04;
input 	mem_95_05;
output 	src_data_95;
input 	mem_96_03;
input 	mem_96_04;
input 	mem_96_05;
output 	src_data_96;
input 	mem_97_03;
input 	mem_97_04;
input 	mem_97_05;
output 	src_data_97;
input 	mem_98_03;
input 	mem_98_04;
input 	mem_98_05;
output 	src_data_98;
input 	mem_99_03;
input 	mem_99_04;
input 	mem_99_05;
output 	src_data_99;
input 	mem_100_03;
input 	mem_100_04;
input 	mem_100_05;
output 	src_data_100;
input 	mem_101_03;
input 	mem_101_04;
input 	mem_101_05;
output 	src_data_101;
input 	mem_102_03;
input 	mem_102_04;
input 	mem_102_05;
output 	src_data_102;
input 	mem_103_03;
input 	mem_103_04;
input 	mem_103_05;
output 	src_data_103;
output 	src_payload22;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~0_combout ;
wire \src_payload~1_combout ;
wire \src_payload~2_combout ;
wire \src_payload~3_combout ;
wire \src_payload~4_combout ;
wire \src_payload~5_combout ;
wire \src_data[0]~0_combout ;
wire \src_data[0]~1_combout ;
wire \src_data[0]~2_combout ;
wire \src_data[0]~3_combout ;
wire \src_data[0]~4_combout ;
wire \src_data[1]~6_combout ;
wire \src_data[1]~7_combout ;
wire \src_data[1]~8_combout ;
wire \src_data[1]~9_combout ;
wire \src_data[1]~10_combout ;
wire \src_data[2]~12_combout ;
wire \src_data[2]~13_combout ;
wire \src_data[2]~14_combout ;
wire \src_payload~6_combout ;
wire \src_data[2]~15_combout ;
wire \src_data[2]~16_combout ;
wire \src_data[3]~18_combout ;
wire \src_data[3]~19_combout ;
wire \src_data[3]~20_combout ;
wire \src_data[3]~21_combout ;
wire \src_data[3]~22_combout ;
wire \src_data[4]~24_combout ;
wire \src_data[4]~25_combout ;
wire \src_data[4]~26_combout ;
wire \src_data[4]~27_combout ;
wire \src_data[4]~28_combout ;
wire \src_data[5]~30_combout ;
wire \src_data[5]~31_combout ;
wire \src_data[5]~32_combout ;
wire \src_data[5]~33_combout ;
wire \src_data[5]~34_combout ;
wire \src_data[6]~36_combout ;
wire \src_data[6]~37_combout ;
wire \src_data[6]~38_combout ;
wire \src_data[6]~39_combout ;
wire \src_data[6]~40_combout ;
wire \src_data[7]~42_combout ;
wire \src_data[7]~43_combout ;
wire \src_data[7]~44_combout ;
wire \src_data[7]~45_combout ;
wire \src_data[7]~46_combout ;
wire \src_data[7]~47_combout ;
wire \src_data[8]~49_combout ;
wire \src_data[8]~50_combout ;
wire \src_data[8]~51_combout ;
wire \src_data[8]~52_combout ;
wire \src_data[8]~53_combout ;
wire \src_payload~7_combout ;
wire \src_data[9]~55_combout ;
wire \src_data[9]~56_combout ;
wire \src_data[9]~57_combout ;
wire \src_data[9]~83_combout ;
wire \src_payload~8_combout ;
wire \src_payload~9_combout ;
wire \src_payload~10_combout ;
wire \src_payload~12_combout ;
wire \src_payload~13_combout ;
wire \src_payload~15_combout ;
wire \src_payload~16_combout ;
wire \src_payload~18_combout ;
wire \src_payload~19_combout ;
wire \src_payload~21_combout ;
wire \src_payload~22_combout ;
wire \src_payload~24_combout ;
wire \src_payload~25_combout ;
wire \src_payload~27_combout ;
wire \src_payload~28_combout ;
wire \src_payload~30_combout ;
wire \src_payload~31_combout ;
wire \src_payload~33_combout ;
wire \src_payload~34_combout ;
wire \src_payload~36_combout ;
wire \src_payload~37_combout ;
wire \src_payload~39_combout ;
wire \src_payload~40_combout ;
wire \src_payload~42_combout ;
wire \src_payload~43_combout ;
wire \src_payload~45_combout ;
wire \src_payload~46_combout ;
wire \src_payload~48_combout ;
wire \src_payload~49_combout ;
wire \src_payload~51_combout ;
wire \src_payload~52_combout ;
wire \src_payload~54_combout ;
wire \src_payload~55_combout ;
wire \src_payload~57_combout ;
wire \src_payload~58_combout ;
wire \src_payload~60_combout ;
wire \src_payload~61_combout ;
wire \src_payload~63_combout ;
wire \src_payload~64_combout ;
wire \src_payload~66_combout ;
wire \src_payload~67_combout ;
wire \src_payload~69_combout ;
wire \src_payload~70_combout ;
wire \src_payload~72_combout ;
wire \src_payload~73_combout ;
wire \src_data[92]~59_combout ;
wire \src_data[92]~60_combout ;
wire \src_data[93]~61_combout ;
wire \src_data[93]~62_combout ;
wire \src_data[94]~63_combout ;
wire \src_data[94]~64_combout ;
wire \src_data[95]~65_combout ;
wire \src_data[95]~66_combout ;
wire \src_data[96]~67_combout ;
wire \src_data[96]~68_combout ;
wire \src_data[97]~69_combout ;
wire \src_data[97]~70_combout ;
wire \src_data[98]~71_combout ;
wire \src_data[98]~72_combout ;
wire \src_data[99]~73_combout ;
wire \src_data[99]~74_combout ;
wire \src_data[100]~75_combout ;
wire \src_data[100]~76_combout ;
wire \src_data[101]~77_combout ;
wire \src_data[101]~78_combout ;
wire \src_data[102]~79_combout ;
wire \src_data[102]~80_combout ;
wire \src_data[103]~81_combout ;
wire \src_data[103]~82_combout ;


cyclonev_lcell_comb \src_payload[0] (
	.dataa(!\src_payload~0_combout ),
	.datab(!\src_payload~1_combout ),
	.datac(!\src_payload~2_combout ),
	.datad(!\src_payload~3_combout ),
	.datae(!\src_payload~4_combout ),
	.dataf(!\src_payload~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload[0] .extended_lut = "off";
defparam \src_payload[0] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload[0] .shared_arith = "off";

cyclonev_lcell_comb WideOr1(
	.dataa(!empty2),
	.datab(!empty1),
	.datac(!empty),
	.datad(!src1_valid),
	.datae(!src1_valid1),
	.dataf(!src1_valid2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~5 (
	.dataa(!\src_data[0]~0_combout ),
	.datab(!\src_data[0]~1_combout ),
	.datac(!\src_data[0]~2_combout ),
	.datad(!\src_data[0]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~5 .extended_lut = "off";
defparam \src_data[0]~5 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~11 (
	.dataa(!\src_data[1]~6_combout ),
	.datab(!\src_data[1]~7_combout ),
	.datac(!\src_data[1]~8_combout ),
	.datad(!\src_data[1]~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~11 .extended_lut = "off";
defparam \src_data[1]~11 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[1]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~17 (
	.dataa(!\src_data[2]~12_combout ),
	.datab(!\src_data[2]~13_combout ),
	.datac(!\src_data[2]~14_combout ),
	.datad(!\src_data[2]~16_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~17 .extended_lut = "off";
defparam \src_data[2]~17 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[2]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~23 (
	.dataa(!\src_data[3]~18_combout ),
	.datab(!\src_data[3]~19_combout ),
	.datac(!\src_data[3]~20_combout ),
	.datad(!\src_data[3]~22_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~23 .extended_lut = "off";
defparam \src_data[3]~23 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[3]~23 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~29 (
	.dataa(!\src_data[4]~24_combout ),
	.datab(!\src_data[4]~25_combout ),
	.datac(!\src_data[4]~26_combout ),
	.datad(!\src_data[4]~28_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~29 .extended_lut = "off";
defparam \src_data[4]~29 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[4]~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~35 (
	.dataa(!\src_data[5]~30_combout ),
	.datab(!\src_data[5]~31_combout ),
	.datac(!\src_data[5]~32_combout ),
	.datad(!\src_data[5]~34_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~35 .extended_lut = "off";
defparam \src_data[5]~35 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[5]~35 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~41 (
	.dataa(!\src_data[6]~36_combout ),
	.datab(!\src_data[6]~37_combout ),
	.datac(!\src_data[6]~38_combout ),
	.datad(!\src_data[6]~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~41 .extended_lut = "off";
defparam \src_data[6]~41 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[6]~41 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~48 (
	.dataa(!\src_data[7]~42_combout ),
	.datab(!\src_data[7]~43_combout ),
	.datac(!\src_data[7]~44_combout ),
	.datad(!\src_data[7]~47_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~48 .extended_lut = "off";
defparam \src_data[7]~48 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[7]~48 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~54 (
	.dataa(!\src_data[8]~49_combout ),
	.datab(!\src_data[8]~50_combout ),
	.datac(!\src_data[8]~51_combout ),
	.datad(!\src_data[8]~53_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~54 .extended_lut = "off";
defparam \src_data[8]~54 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src_data[8]~54 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~58 (
	.dataa(!\src_payload~7_combout ),
	.datab(!\src_data[9]~55_combout ),
	.datac(!\src_data[9]~56_combout ),
	.datad(!\src_data[9]~57_combout ),
	.datae(!\src_data[9]~83_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~58 .extended_lut = "off";
defparam \src_data[9]~58 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[9]~58 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!\src_data[7]~45_combout ),
	.datab(!\src_payload~8_combout ),
	.datac(!\src_payload~9_combout ),
	.datad(!\src_payload~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_111),
	.datad(!mem_11_01),
	.datae(!\src_payload~12_combout ),
	.dataf(!\src_payload~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_121),
	.datad(!mem_12_0),
	.datae(!\src_payload~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_131),
	.datad(!mem_13_0),
	.datae(!\src_payload~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_141),
	.datad(!mem_14_0),
	.datae(!\src_payload~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_15),
	.datad(!mem_15_0),
	.datae(!\src_payload~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_16),
	.datad(!mem_16_0),
	.datae(!\src_payload~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_17),
	.datad(!mem_17_0),
	.datae(!\src_payload~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~35 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_18),
	.datad(!mem_18_0),
	.datae(!\src_payload~34_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~35 .extended_lut = "off";
defparam \src_payload~35 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~35 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~38 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_19),
	.datad(!mem_19_0),
	.datae(!\src_payload~36_combout ),
	.dataf(!\src_payload~37_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~38 .extended_lut = "off";
defparam \src_payload~38 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~38 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~41 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_20),
	.datad(!mem_20_0),
	.datae(!\src_payload~39_combout ),
	.dataf(!\src_payload~40_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~41 .extended_lut = "off";
defparam \src_payload~41 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~41 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~44 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_211),
	.datad(!mem_21_0),
	.datae(!\src_payload~42_combout ),
	.dataf(!\src_payload~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~44 .extended_lut = "off";
defparam \src_payload~44 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~44 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~47 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_221),
	.datad(!mem_22_0),
	.datae(!\src_payload~46_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~47 .extended_lut = "off";
defparam \src_payload~47 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~47 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~50 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_231),
	.datad(!mem_23_0),
	.datae(!\src_payload~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~50 .extended_lut = "off";
defparam \src_payload~50 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~50 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~53 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_241),
	.datad(!mem_24_0),
	.datae(!\src_payload~51_combout ),
	.dataf(!\src_payload~52_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~53 .extended_lut = "off";
defparam \src_payload~53 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~53 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~56 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_25),
	.datad(!mem_25_0),
	.datae(!\src_payload~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~56 .extended_lut = "off";
defparam \src_payload~56 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~56 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~59 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_26),
	.datad(!mem_26_0),
	.datae(!\src_payload~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~59 .extended_lut = "off";
defparam \src_payload~59 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~59 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~62 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_27),
	.datad(!mem_27_0),
	.datae(!\src_payload~60_combout ),
	.dataf(!\src_payload~61_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~62 .extended_lut = "off";
defparam \src_payload~62 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~62 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~65 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_28),
	.datad(!mem_28_0),
	.datae(!\src_payload~63_combout ),
	.dataf(!\src_payload~64_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~65 .extended_lut = "off";
defparam \src_payload~65 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~65 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~68 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_29),
	.datad(!mem_29_0),
	.datae(!\src_payload~67_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~68 .extended_lut = "off";
defparam \src_payload~68 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~68 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~71 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_301),
	.datad(!mem_30_0),
	.datae(!\src_payload~69_combout ),
	.dataf(!\src_payload~70_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~71 .extended_lut = "off";
defparam \src_payload~71 .lut_mask = 64'hFFFFFFFF028AFFFF;
defparam \src_payload~71 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~74 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_311),
	.datad(!mem_31_0),
	.datae(!\src_payload~73_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~74 .extended_lut = "off";
defparam \src_payload~74 .lut_mask = 64'hFFFF028AFFFF028A;
defparam \src_payload~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_92_01),
	.datad(!mem_92_02),
	.datae(!\src_data[92]~60_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_92),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92] .extended_lut = "off";
defparam \src_data[92] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[92] .shared_arith = "off";

cyclonev_lcell_comb \src_data[93] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_93_01),
	.datad(!mem_93_02),
	.datae(!\src_data[93]~62_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_93),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93] .extended_lut = "off";
defparam \src_data[93] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[93] .shared_arith = "off";

cyclonev_lcell_comb \src_data[94] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_94_01),
	.datad(!mem_94_02),
	.datae(!\src_data[94]~64_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_94),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94] .extended_lut = "off";
defparam \src_data[94] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[94] .shared_arith = "off";

cyclonev_lcell_comb \src_data[95] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_95_01),
	.datad(!mem_95_02),
	.datae(!\src_data[95]~66_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_95),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95] .extended_lut = "off";
defparam \src_data[95] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[95] .shared_arith = "off";

cyclonev_lcell_comb \src_data[96] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_96_01),
	.datad(!mem_96_02),
	.datae(!\src_data[96]~68_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_96),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96] .extended_lut = "off";
defparam \src_data[96] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[96] .shared_arith = "off";

cyclonev_lcell_comb \src_data[97] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_97_01),
	.datad(!mem_97_02),
	.datae(!\src_data[97]~70_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_97),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97] .extended_lut = "off";
defparam \src_data[97] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[97] .shared_arith = "off";

cyclonev_lcell_comb \src_data[98] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_98_01),
	.datad(!mem_98_02),
	.datae(!\src_data[98]~72_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_98),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98] .extended_lut = "off";
defparam \src_data[98] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[98] .shared_arith = "off";

cyclonev_lcell_comb \src_data[99] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_99_01),
	.datad(!mem_99_02),
	.datae(!\src_data[99]~74_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_99),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99] .extended_lut = "off";
defparam \src_data[99] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[99] .shared_arith = "off";

cyclonev_lcell_comb \src_data[100] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_100_01),
	.datad(!mem_100_02),
	.datae(!\src_data[100]~76_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_100),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100] .extended_lut = "off";
defparam \src_data[100] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[100] .shared_arith = "off";

cyclonev_lcell_comb \src_data[101] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_101_01),
	.datad(!mem_101_02),
	.datae(!\src_data[101]~78_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_101),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101] .extended_lut = "off";
defparam \src_data[101] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[101] .shared_arith = "off";

cyclonev_lcell_comb \src_data[102] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_102_01),
	.datad(!mem_102_02),
	.datae(!\src_data[102]~80_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_102),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102] .extended_lut = "off";
defparam \src_data[102] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[102] .shared_arith = "off";

cyclonev_lcell_comb \src_data[103] (
	.dataa(!src1_valid1),
	.datab(!src1_valid2),
	.datac(!mem_103_01),
	.datad(!mem_103_02),
	.datae(!\src_data[103]~82_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_103),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103] .extended_lut = "off";
defparam \src_data[103] .lut_mask = 64'hFFFF0ACEFFFF0ACE;
defparam \src_data[103] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~75 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!mem_117_0),
	.datad(!last_packet_beat),
	.datae(!last_packet_beat1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~75 .extended_lut = "off";
defparam \src_payload~75 .lut_mask = 64'h0C0D0D0D0C0D0D0D;
defparam \src_payload~75 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!comb),
	.datab(!mem_57_0),
	.datac(!src1_valid),
	.datad(!mem_117_0),
	.datae(!last_packet_beat),
	.dataf(!last_packet_beat1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!comb1),
	.datab(!mem_57_01),
	.datac(!src1_valid1),
	.datad(!mem_117_01),
	.datae(!last_packet_beat2),
	.dataf(!last_packet_beat3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!comb2),
	.datab(!mem_57_02),
	.datac(!src1_valid2),
	.datad(!mem_117_02),
	.datae(!last_packet_beat4),
	.dataf(!last_packet_beat5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h00C000D000D000D0;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!mem_117_03),
	.datab(!empty),
	.datac(!mem_57_03),
	.datad(!mem_used_01),
	.datae(!last_packet_beat6),
	.dataf(!last_packet_beat7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h4040404440444044;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!mem_117_04),
	.datab(!empty1),
	.datac(!mem_57_04),
	.datad(!mem_used_03),
	.datae(!last_packet_beat8),
	.dataf(!last_packet_beat9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h4040404440444044;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!mem_117_05),
	.datab(!empty2),
	.datac(!mem_57_05),
	.datad(!mem_used_05),
	.datae(!last_packet_beat10),
	.dataf(!last_packet_beat11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h4040404440444044;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!src1_valid),
	.datab(!av_readdata_pre_0),
	.datac(!always4),
	.datad(!mem_0_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'h02A202A202A202A2;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!src1_valid1),
	.datab(!av_readdata_pre_01),
	.datac(!always41),
	.datad(!mem_0_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'h02A202A202A202A2;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~2 (
	.dataa(!src1_valid2),
	.datab(!av_readdata_pre_02),
	.datac(!always42),
	.datad(!mem_0_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~2 .extended_lut = "off";
defparam \src_data[0]~2 .lut_mask = 64'h02A202A202A202A2;
defparam \src_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_0_04),
	.datad(!av_readdata_pre_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~3 .extended_lut = "off";
defparam \src_data[0]~3 .lut_mask = 64'h0347034703470347;
defparam \src_data[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~4 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_0_03),
	.datad(!av_readdata_pre_03),
	.datae(!\src_data[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~4 .extended_lut = "off";
defparam \src_data[0]~4 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[0]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~6 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_1),
	.datad(!mem_1_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~6 .extended_lut = "off";
defparam \src_data[1]~6 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~7 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_11),
	.datad(!mem_1_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~7 .extended_lut = "off";
defparam \src_data[1]~7 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~8 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_12),
	.datad(!mem_1_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~8 .extended_lut = "off";
defparam \src_data[1]~8 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[1]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~9 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_1_04),
	.datad(!av_readdata_pre_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~9 .extended_lut = "off";
defparam \src_data[1]~9 .lut_mask = 64'h0347034703470347;
defparam \src_data[1]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~10 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_1_03),
	.datad(!av_readdata_pre_13),
	.datae(!\src_data[1]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~10 .extended_lut = "off";
defparam \src_data[1]~10 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[1]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~12 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_2),
	.datad(!mem_2_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~12 .extended_lut = "off";
defparam \src_data[2]~12 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[2]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~13 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_21),
	.datad(!mem_2_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~13 .extended_lut = "off";
defparam \src_data[2]~13 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[2]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~14 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_22),
	.datad(!mem_2_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~14 .extended_lut = "off";
defparam \src_data[2]~14 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[2]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!mem_11_0),
	.datad(!av_readdata_pre_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h0347034703470347;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~15 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_2_04),
	.datad(!av_readdata_pre_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~15 .extended_lut = "off";
defparam \src_data[2]~15 .lut_mask = 64'h0347034703470347;
defparam \src_data[2]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~16 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_2_03),
	.datad(!av_readdata_pre_23),
	.datae(!\src_payload~6_combout ),
	.dataf(!\src_data[2]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~16 .extended_lut = "off";
defparam \src_data[2]~16 .lut_mask = 64'hFCB8000000000000;
defparam \src_data[2]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~18 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_3),
	.datad(!mem_3_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~18 .extended_lut = "off";
defparam \src_data[3]~18 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[3]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~19 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_31),
	.datad(!mem_3_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~19 .extended_lut = "off";
defparam \src_data[3]~19 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[3]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~20 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_32),
	.datad(!mem_3_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~20 .extended_lut = "off";
defparam \src_data[3]~20 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[3]~20 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~21 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_3_04),
	.datad(!av_readdata_pre_34),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~21 .extended_lut = "off";
defparam \src_data[3]~21 .lut_mask = 64'h0347034703470347;
defparam \src_data[3]~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~22 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_3_03),
	.datad(!av_readdata_pre_33),
	.datae(!\src_data[3]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~22 .extended_lut = "off";
defparam \src_data[3]~22 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[3]~22 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~24 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_4),
	.datad(!mem_4_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~24 .extended_lut = "off";
defparam \src_data[4]~24 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[4]~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~25 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_41),
	.datad(!mem_4_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~25 .extended_lut = "off";
defparam \src_data[4]~25 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[4]~25 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~26 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_42),
	.datad(!mem_4_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~26 .extended_lut = "off";
defparam \src_data[4]~26 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[4]~26 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~27 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_4_04),
	.datad(!av_readdata_pre_44),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~27 .extended_lut = "off";
defparam \src_data[4]~27 .lut_mask = 64'h0347034703470347;
defparam \src_data[4]~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~28 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_4_03),
	.datad(!av_readdata_pre_43),
	.datae(!\src_data[4]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~28 .extended_lut = "off";
defparam \src_data[4]~28 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[4]~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~30 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_5),
	.datad(!mem_5_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~30 .extended_lut = "off";
defparam \src_data[5]~30 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[5]~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~31 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_51),
	.datad(!mem_5_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~31 .extended_lut = "off";
defparam \src_data[5]~31 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[5]~31 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~32 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_52),
	.datad(!mem_5_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~32 .extended_lut = "off";
defparam \src_data[5]~32 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[5]~32 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~33 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_5_04),
	.datad(!av_readdata_pre_54),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~33 .extended_lut = "off";
defparam \src_data[5]~33 .lut_mask = 64'h0347034703470347;
defparam \src_data[5]~33 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~34 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_5_03),
	.datad(!av_readdata_pre_53),
	.datae(!\src_data[5]~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~34 .extended_lut = "off";
defparam \src_data[5]~34 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[5]~34 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~36 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_6),
	.datad(!mem_6_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~36 .extended_lut = "off";
defparam \src_data[6]~36 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[6]~36 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~37 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_61),
	.datad(!mem_6_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~37 .extended_lut = "off";
defparam \src_data[6]~37 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[6]~37 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~38 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_62),
	.datad(!mem_6_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~38 .extended_lut = "off";
defparam \src_data[6]~38 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[6]~38 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~39 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_6_04),
	.datad(!av_readdata_pre_64),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~39 .extended_lut = "off";
defparam \src_data[6]~39 .lut_mask = 64'h0347034703470347;
defparam \src_data[6]~39 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~40 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_6_03),
	.datad(!av_readdata_pre_63),
	.datae(!\src_data[6]~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~40 .extended_lut = "off";
defparam \src_data[6]~40 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[6]~40 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~42 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_7),
	.datad(!mem_7_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~42 .extended_lut = "off";
defparam \src_data[7]~42 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[7]~42 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~43 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_71),
	.datad(!mem_7_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~43 .extended_lut = "off";
defparam \src_data[7]~43 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[7]~43 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~44 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_72),
	.datad(!mem_7_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~44 .extended_lut = "off";
defparam \src_data[7]~44 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[7]~44 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~45 (
	.dataa(!in_ready_hold),
	.datab(!read_latency_shift_reg_02),
	.datac(!mem_used_04),
	.datad(!mem_10_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~45 .extended_lut = "off";
defparam \src_data[7]~45 .lut_mask = 64'h101F101F101F101F;
defparam \src_data[7]~45 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~46 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_7_04),
	.datad(!av_readdata_pre_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~46 .extended_lut = "off";
defparam \src_data[7]~46 .lut_mask = 64'h0347034703470347;
defparam \src_data[7]~46 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~47 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_7_03),
	.datad(!av_readdata_pre_73),
	.datae(!\src_data[7]~45_combout ),
	.dataf(!\src_data[7]~46_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~47 .extended_lut = "off";
defparam \src_data[7]~47 .lut_mask = 64'hFCB8000000000000;
defparam \src_data[7]~47 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~49 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_8),
	.datad(!mem_8_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~49 .extended_lut = "off";
defparam \src_data[8]~49 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[8]~49 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~50 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_81),
	.datad(!mem_8_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~50 .extended_lut = "off";
defparam \src_data[8]~50 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[8]~50 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~51 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_82),
	.datad(!mem_8_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~51 .extended_lut = "off";
defparam \src_data[8]~51 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[8]~51 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~52 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_0),
	.datac(!mem_8_04),
	.datad(!av_readdata_pre_84),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~52 .extended_lut = "off";
defparam \src_data[8]~52 .lut_mask = 64'h0347034703470347;
defparam \src_data[8]~52 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~53 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_8_03),
	.datad(!av_readdata_pre_83),
	.datae(!\src_data[8]~52_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~53 .extended_lut = "off";
defparam \src_data[8]~53 .lut_mask = 64'hFCB80000FCB80000;
defparam \src_data[8]~53 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!av_readdata_pre_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h0404040404040404;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~55 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_91),
	.datad(!mem_9_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~55 .extended_lut = "off";
defparam \src_data[9]~55 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[9]~55 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~56 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_92),
	.datad(!mem_9_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~56 .extended_lut = "off";
defparam \src_data[9]~56 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[9]~56 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~57 (
	.dataa(!src1_valid2),
	.datab(!always42),
	.datac(!av_readdata_pre_93),
	.datad(!mem_9_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~57 .extended_lut = "off";
defparam \src_data[9]~57 .lut_mask = 64'h028A028A028A028A;
defparam \src_data[9]~57 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~83 (
	.dataa(!mem_9_04),
	.datab(!av_readdata_pre_94),
	.datac(!mem_9_03),
	.datad(!mem_used_02),
	.datae(!mem_used_0),
	.dataf(!\src_payload~6_combout ),
	.datag(!read_latency_shift_reg_0),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~83 .extended_lut = "on";
defparam \src_data[9]~83 .lut_mask = 64'h03570F5FFFFFFFFF;
defparam \src_data[9]~83 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_10),
	.datad(!mem_10_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_101),
	.datad(!mem_10_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_10_03),
	.datad(!av_readdata_pre_102),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h0347034703470347;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_112),
	.datad(!mem_11_02),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_11_03),
	.datae(!av_readdata_pre_113),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_12_02),
	.datad(!av_readdata_pre_123),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h0347034703470347;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_122),
	.datad(!mem_12_01),
	.datae(!\src_payload~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_13_02),
	.datad(!av_readdata_pre_133),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h0347034703470347;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_132),
	.datad(!mem_13_01),
	.datae(!\src_payload~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_14_02),
	.datad(!av_readdata_pre_143),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h0347034703470347;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_142),
	.datad(!mem_14_01),
	.datae(!\src_payload~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_15_02),
	.datad(!av_readdata_pre_152),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h0347034703470347;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_151),
	.datad(!mem_15_01),
	.datae(!\src_payload~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_16_02),
	.datad(!av_readdata_pre_162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h0347034703470347;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_161),
	.datad(!mem_16_01),
	.datae(!\src_payload~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_17_02),
	.datad(!av_readdata_pre_172),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h0347034703470347;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_171),
	.datad(!mem_17_01),
	.datae(!\src_payload~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~33 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_18_02),
	.datad(!av_readdata_pre_182),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~33 .extended_lut = "off";
defparam \src_payload~33 .lut_mask = 64'h0347034703470347;
defparam \src_payload~33 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~34 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_181),
	.datad(!mem_18_01),
	.datae(!\src_payload~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~34 .extended_lut = "off";
defparam \src_payload~34 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~34 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~36 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_191),
	.datad(!mem_19_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~36 .extended_lut = "off";
defparam \src_payload~36 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~36 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~37 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_19_02),
	.datae(!av_readdata_pre_192),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~37 .extended_lut = "off";
defparam \src_payload~37 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~37 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~39 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_201),
	.datad(!mem_20_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~39 .extended_lut = "off";
defparam \src_payload~39 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~39 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~40 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_20_02),
	.datae(!av_readdata_pre_202),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~40 .extended_lut = "off";
defparam \src_payload~40 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~40 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~42 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_212),
	.datad(!mem_21_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~42 .extended_lut = "off";
defparam \src_payload~42 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~42 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~43 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_21_02),
	.datae(!av_readdata_pre_213),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~43 .extended_lut = "off";
defparam \src_payload~43 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~43 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~45 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_22_02),
	.datad(!av_readdata_pre_223),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~45 .extended_lut = "off";
defparam \src_payload~45 .lut_mask = 64'h0347034703470347;
defparam \src_payload~45 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~46 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_222),
	.datad(!mem_22_01),
	.datae(!\src_payload~45_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~46 .extended_lut = "off";
defparam \src_payload~46 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~46 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~48 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_23_02),
	.datad(!av_readdata_pre_233),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~48 .extended_lut = "off";
defparam \src_payload~48 .lut_mask = 64'h0347034703470347;
defparam \src_payload~48 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~49 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_232),
	.datad(!mem_23_01),
	.datae(!\src_payload~48_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~49 .extended_lut = "off";
defparam \src_payload~49 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~49 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~51 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_242),
	.datad(!mem_24_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~51 .extended_lut = "off";
defparam \src_payload~51 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~51 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~52 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_24_02),
	.datae(!av_readdata_pre_243),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~52 .extended_lut = "off";
defparam \src_payload~52 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~52 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~54 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_25_02),
	.datad(!av_readdata_pre_252),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~54 .extended_lut = "off";
defparam \src_payload~54 .lut_mask = 64'h0347034703470347;
defparam \src_payload~54 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~55 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_251),
	.datad(!mem_25_01),
	.datae(!\src_payload~54_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~55 .extended_lut = "off";
defparam \src_payload~55 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~55 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~57 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_26_02),
	.datad(!av_readdata_pre_262),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~57 .extended_lut = "off";
defparam \src_payload~57 .lut_mask = 64'h0347034703470347;
defparam \src_payload~57 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~58 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_261),
	.datad(!mem_26_01),
	.datae(!\src_payload~57_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~58 .extended_lut = "off";
defparam \src_payload~58 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~58 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~60 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_271),
	.datad(!mem_27_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~60 .extended_lut = "off";
defparam \src_payload~60 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~60 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~61 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_27_02),
	.datae(!av_readdata_pre_272),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~61 .extended_lut = "off";
defparam \src_payload~61 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~61 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~63 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_281),
	.datad(!mem_28_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~63 .extended_lut = "off";
defparam \src_payload~63 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~63 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~64 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_28_02),
	.datae(!av_readdata_pre_282),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~64 .extended_lut = "off";
defparam \src_payload~64 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~64 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~66 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_29_02),
	.datad(!av_readdata_pre_292),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~66 .extended_lut = "off";
defparam \src_payload~66 .lut_mask = 64'h0347034703470347;
defparam \src_payload~66 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~67 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_291),
	.datad(!mem_29_01),
	.datae(!\src_payload~66_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~67 .extended_lut = "off";
defparam \src_payload~67 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~67 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~69 (
	.dataa(!src1_valid1),
	.datab(!always41),
	.datac(!av_readdata_pre_302),
	.datad(!mem_30_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~69 .extended_lut = "off";
defparam \src_payload~69 .lut_mask = 64'h028A028A028A028A;
defparam \src_payload~69 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~70 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!\src_payload~6_combout ),
	.datad(!mem_30_02),
	.datae(!av_readdata_pre_303),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~70 .extended_lut = "off";
defparam \src_payload~70 .lut_mask = 64'hF0C0B080F0C0B080;
defparam \src_payload~70 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~72 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!mem_used_02),
	.datac(!mem_31_02),
	.datad(!av_readdata_pre_313),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~72 .extended_lut = "off";
defparam \src_payload~72 .lut_mask = 64'h0347034703470347;
defparam \src_payload~72 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~73 (
	.dataa(!src1_valid),
	.datab(!always4),
	.datac(!av_readdata_pre_312),
	.datad(!mem_31_01),
	.datae(!\src_payload~72_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~73 .extended_lut = "off";
defparam \src_payload~73 .lut_mask = 64'hFD750000FD750000;
defparam \src_payload~73 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92]~59 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_92_04),
	.dataf(!mem_92_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[92]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92]~59 .extended_lut = "off";
defparam \src_data[92]~59 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[92]~59 .shared_arith = "off";

cyclonev_lcell_comb \src_data[92]~60 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_92_0),
	.datad(!mem_92_03),
	.datae(!\src_data[92]~59_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[92]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[92]~60 .extended_lut = "off";
defparam \src_data[92]~60 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[92]~60 .shared_arith = "off";

cyclonev_lcell_comb \src_data[93]~61 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_93_04),
	.dataf(!mem_93_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[93]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93]~61 .extended_lut = "off";
defparam \src_data[93]~61 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[93]~61 .shared_arith = "off";

cyclonev_lcell_comb \src_data[93]~62 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_93_0),
	.datad(!mem_93_03),
	.datae(!\src_data[93]~61_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[93]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[93]~62 .extended_lut = "off";
defparam \src_data[93]~62 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[93]~62 .shared_arith = "off";

cyclonev_lcell_comb \src_data[94]~63 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_94_04),
	.dataf(!mem_94_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[94]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94]~63 .extended_lut = "off";
defparam \src_data[94]~63 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[94]~63 .shared_arith = "off";

cyclonev_lcell_comb \src_data[94]~64 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_94_0),
	.datad(!mem_94_03),
	.datae(!\src_data[94]~63_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[94]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[94]~64 .extended_lut = "off";
defparam \src_data[94]~64 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[94]~64 .shared_arith = "off";

cyclonev_lcell_comb \src_data[95]~65 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_95_04),
	.dataf(!mem_95_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[95]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95]~65 .extended_lut = "off";
defparam \src_data[95]~65 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[95]~65 .shared_arith = "off";

cyclonev_lcell_comb \src_data[95]~66 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_95_0),
	.datad(!mem_95_03),
	.datae(!\src_data[95]~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[95]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[95]~66 .extended_lut = "off";
defparam \src_data[95]~66 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[95]~66 .shared_arith = "off";

cyclonev_lcell_comb \src_data[96]~67 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_96_04),
	.dataf(!mem_96_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[96]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96]~67 .extended_lut = "off";
defparam \src_data[96]~67 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[96]~67 .shared_arith = "off";

cyclonev_lcell_comb \src_data[96]~68 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_96_0),
	.datad(!mem_96_03),
	.datae(!\src_data[96]~67_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[96]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[96]~68 .extended_lut = "off";
defparam \src_data[96]~68 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[96]~68 .shared_arith = "off";

cyclonev_lcell_comb \src_data[97]~69 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_97_04),
	.dataf(!mem_97_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[97]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97]~69 .extended_lut = "off";
defparam \src_data[97]~69 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[97]~69 .shared_arith = "off";

cyclonev_lcell_comb \src_data[97]~70 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_97_0),
	.datad(!mem_97_03),
	.datae(!\src_data[97]~69_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[97]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[97]~70 .extended_lut = "off";
defparam \src_data[97]~70 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[97]~70 .shared_arith = "off";

cyclonev_lcell_comb \src_data[98]~71 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_98_04),
	.dataf(!mem_98_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[98]~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98]~71 .extended_lut = "off";
defparam \src_data[98]~71 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[98]~71 .shared_arith = "off";

cyclonev_lcell_comb \src_data[98]~72 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_98_0),
	.datad(!mem_98_03),
	.datae(!\src_data[98]~71_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[98]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[98]~72 .extended_lut = "off";
defparam \src_data[98]~72 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[98]~72 .shared_arith = "off";

cyclonev_lcell_comb \src_data[99]~73 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_99_04),
	.dataf(!mem_99_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[99]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99]~73 .extended_lut = "off";
defparam \src_data[99]~73 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[99]~73 .shared_arith = "off";

cyclonev_lcell_comb \src_data[99]~74 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_99_0),
	.datad(!mem_99_03),
	.datae(!\src_data[99]~73_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[99]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[99]~74 .extended_lut = "off";
defparam \src_data[99]~74 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[99]~74 .shared_arith = "off";

cyclonev_lcell_comb \src_data[100]~75 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_100_04),
	.dataf(!mem_100_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[100]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100]~75 .extended_lut = "off";
defparam \src_data[100]~75 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[100]~75 .shared_arith = "off";

cyclonev_lcell_comb \src_data[100]~76 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_100_0),
	.datad(!mem_100_03),
	.datae(!\src_data[100]~75_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[100]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[100]~76 .extended_lut = "off";
defparam \src_data[100]~76 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[100]~76 .shared_arith = "off";

cyclonev_lcell_comb \src_data[101]~77 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_101_04),
	.dataf(!mem_101_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[101]~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101]~77 .extended_lut = "off";
defparam \src_data[101]~77 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[101]~77 .shared_arith = "off";

cyclonev_lcell_comb \src_data[101]~78 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_101_0),
	.datad(!mem_101_03),
	.datae(!\src_data[101]~77_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[101]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[101]~78 .extended_lut = "off";
defparam \src_data[101]~78 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[101]~78 .shared_arith = "off";

cyclonev_lcell_comb \src_data[102]~79 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_102_04),
	.dataf(!mem_102_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[102]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102]~79 .extended_lut = "off";
defparam \src_data[102]~79 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[102]~79 .shared_arith = "off";

cyclonev_lcell_comb \src_data[102]~80 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_102_0),
	.datad(!mem_102_03),
	.datae(!\src_data[102]~79_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[102]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[102]~80 .extended_lut = "off";
defparam \src_data[102]~80 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[102]~80 .shared_arith = "off";

cyclonev_lcell_comb \src_data[103]~81 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!mem_used_04),
	.datac(!read_latency_shift_reg_01),
	.datad(!mem_used_02),
	.datae(!mem_103_04),
	.dataf(!mem_103_05),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[103]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103]~81 .extended_lut = "off";
defparam \src_data[103]~81 .lut_mask = 64'hFFFF8888F0008000;
defparam \src_data[103]~81 .shared_arith = "off";

cyclonev_lcell_comb \src_data[103]~82 (
	.dataa(!empty),
	.datab(!src1_valid),
	.datac(!mem_103_0),
	.datad(!mem_103_03),
	.datae(!\src_data[103]~81_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[103]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[103]~82 .extended_lut = "off";
defparam \src_data[103]~82 .lut_mask = 64'h0000F3510000F351;
defparam \src_data[103]~82 .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_rst_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_reset_controller_1 rst_controller(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk_clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module terminal_qsys_terminal_qsys_rst_controller_1 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_reset_controller rst_controller(
	.h2f_rst_n_0(h2f_rst_n_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk_clk(clk_clk));

endmodule

module terminal_qsys_altera_reset_controller (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.h2f_rst_n_0(h2f_rst_n_0),
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

endmodule

module terminal_qsys_altera_reset_synchronizer_1 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(h2f_rst_n_0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module terminal_qsys_altera_reset_controller_1 (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module terminal_qsys_altera_reset_synchronizer_3 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module terminal_qsys_terminal_qsys_rst_controller_001 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



terminal_qsys_altera_reset_controller_2 rst_controller_001(
	.h2f_rst_n_0(h2f_rst_n_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk_clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module terminal_qsys_altera_reset_controller_2 (
	h2f_rst_n_0,
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	h2f_rst_n_0;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \merged_reset~0_combout ;


terminal_qsys_altera_reset_synchronizer_5 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.merged_reset(\merged_reset~0_combout ),
	.clk(clk_clk));

cyclonev_lcell_comb \merged_reset~0 (
	.dataa(!h2f_rst_n_0),
	.datab(!reset_reset_n),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\merged_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_reset~0 .extended_lut = "off";
defparam \merged_reset~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \merged_reset~0 .shared_arith = "off";

endmodule

module terminal_qsys_altera_reset_synchronizer_5 (
	altera_reset_synchronizer_int_chain_out1,
	merged_reset,
	clk)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	merged_reset;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!merged_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module terminal_qsys_terminal_qsys_state (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	readdata_10,
	readdata_11,
	readdata_12,
	readdata_13,
	readdata_14,
	readdata_15,
	readdata_16,
	readdata_17,
	readdata_18,
	readdata_19,
	readdata_20,
	readdata_21,
	readdata_22,
	readdata_23,
	readdata_24,
	readdata_25,
	readdata_26,
	readdata_27,
	readdata_28,
	readdata_29,
	readdata_30,
	readdata_31,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	state_in_export_0,
	state_in_export_1,
	state_in_export_2,
	state_in_export_3,
	state_in_export_4,
	state_in_export_5,
	state_in_export_6,
	state_in_export_7,
	state_in_export_8,
	state_in_export_9,
	state_in_export_10,
	state_in_export_11,
	state_in_export_12,
	state_in_export_13,
	state_in_export_14,
	state_in_export_15,
	state_in_export_16,
	state_in_export_17,
	state_in_export_18,
	state_in_export_19,
	state_in_export_20,
	state_in_export_21,
	state_in_export_22,
	state_in_export_23,
	state_in_export_24,
	state_in_export_25,
	state_in_export_26,
	state_in_export_27,
	state_in_export_28,
	state_in_export_29,
	state_in_export_30,
	state_in_export_31)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
output 	readdata_10;
output 	readdata_11;
output 	readdata_12;
output 	readdata_13;
output 	readdata_14;
output 	readdata_15;
output 	readdata_16;
output 	readdata_17;
output 	readdata_18;
output 	readdata_19;
output 	readdata_20;
output 	readdata_21;
output 	readdata_22;
output 	readdata_23;
output 	readdata_24;
output 	readdata_25;
output 	readdata_26;
output 	readdata_27;
output 	readdata_28;
output 	readdata_29;
output 	readdata_30;
output 	readdata_31;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	state_in_export_0;
input 	state_in_export_1;
input 	state_in_export_2;
input 	state_in_export_3;
input 	state_in_export_4;
input 	state_in_export_5;
input 	state_in_export_6;
input 	state_in_export_7;
input 	state_in_export_8;
input 	state_in_export_9;
input 	state_in_export_10;
input 	state_in_export_11;
input 	state_in_export_12;
input 	state_in_export_13;
input 	state_in_export_14;
input 	state_in_export_15;
input 	state_in_export_16;
input 	state_in_export_17;
input 	state_in_export_18;
input 	state_in_export_19;
input 	state_in_export_20;
input 	state_in_export_21;
input 	state_in_export_22;
input 	state_in_export_23;
input 	state_in_export_24;
input 	state_in_export_25;
input 	state_in_export_26;
input 	state_in_export_27;
input 	state_in_export_28;
input 	state_in_export_29;
input 	state_in_export_30;
input 	state_in_export_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;
wire \read_mux_out[8]~combout ;
wire \read_mux_out[9]~combout ;
wire \read_mux_out[10]~combout ;
wire \read_mux_out[11]~combout ;
wire \read_mux_out[12]~combout ;
wire \read_mux_out[13]~combout ;
wire \read_mux_out[14]~combout ;
wire \read_mux_out[15]~combout ;
wire \read_mux_out[16]~combout ;
wire \read_mux_out[17]~combout ;
wire \read_mux_out[18]~combout ;
wire \read_mux_out[19]~combout ;
wire \read_mux_out[20]~combout ;
wire \read_mux_out[21]~combout ;
wire \read_mux_out[22]~combout ;
wire \read_mux_out[23]~combout ;
wire \read_mux_out[24]~combout ;
wire \read_mux_out[25]~combout ;
wire \read_mux_out[26]~combout ;
wire \read_mux_out[27]~combout ;
wire \read_mux_out[28]~combout ;
wire \read_mux_out[29]~combout ;
wire \read_mux_out[30]~combout ;
wire \read_mux_out[31]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\read_mux_out[8]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\read_mux_out[9]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\read_mux_out[10]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\read_mux_out[11]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\read_mux_out[12]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\read_mux_out[13]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\read_mux_out[14]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\read_mux_out[15]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\read_mux_out[16]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\read_mux_out[17]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\read_mux_out[18]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\read_mux_out[19]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\read_mux_out[20]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\read_mux_out[21]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\read_mux_out[22]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\read_mux_out[23]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\read_mux_out[24]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\read_mux_out[25]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\read_mux_out[26]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\read_mux_out[27]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\read_mux_out[28]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\read_mux_out[29]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\read_mux_out[30]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\read_mux_out[31]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!state_in_export_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h4040404040404040;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[7] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[8] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8] .extended_lut = "off";
defparam \read_mux_out[8] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[8] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[9] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[9] .extended_lut = "off";
defparam \read_mux_out[9] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[9] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[10] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[10] .extended_lut = "off";
defparam \read_mux_out[10] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[10] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[11] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[11] .extended_lut = "off";
defparam \read_mux_out[11] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[11] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[12] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[12] .extended_lut = "off";
defparam \read_mux_out[12] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[12] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[13] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[13] .extended_lut = "off";
defparam \read_mux_out[13] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[13] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[14] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[14] .extended_lut = "off";
defparam \read_mux_out[14] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[14] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[15] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[15] .extended_lut = "off";
defparam \read_mux_out[15] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[15] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[16] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[16] .extended_lut = "off";
defparam \read_mux_out[16] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[16] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[17] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[17] .extended_lut = "off";
defparam \read_mux_out[17] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[17] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[18] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[18] .extended_lut = "off";
defparam \read_mux_out[18] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[18] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[19] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[19] .extended_lut = "off";
defparam \read_mux_out[19] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[19] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[20] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[20] .extended_lut = "off";
defparam \read_mux_out[20] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[20] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[21] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[21] .extended_lut = "off";
defparam \read_mux_out[21] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[21] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[22] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[22] .extended_lut = "off";
defparam \read_mux_out[22] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[22] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[23] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[23] .extended_lut = "off";
defparam \read_mux_out[23] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[23] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[24] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[24] .extended_lut = "off";
defparam \read_mux_out[24] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[24] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[25] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[25] .extended_lut = "off";
defparam \read_mux_out[25] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[25] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[26] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[26] .extended_lut = "off";
defparam \read_mux_out[26] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[26] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[27] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[27] .extended_lut = "off";
defparam \read_mux_out[27] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[27] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[28] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[28] .extended_lut = "off";
defparam \read_mux_out[28] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[28] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[29] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[29] .extended_lut = "off";
defparam \read_mux_out[29] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[29] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[30] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[30] .extended_lut = "off";
defparam \read_mux_out[30] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[30] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[31] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!state_in_export_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[31] .extended_lut = "off";
defparam \read_mux_out[31] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[31] .shared_arith = "off";

endmodule

module terminal_qsys_terminal_qsys_switches (
	altera_reset_synchronizer_int_chain_out,
	readdata_0,
	readdata_1,
	readdata_2,
	readdata_3,
	readdata_4,
	readdata_5,
	readdata_6,
	readdata_7,
	readdata_8,
	readdata_9,
	int_nxt_addr_reg_dly_3,
	int_nxt_addr_reg_dly_2,
	clk_clk,
	switches_in_export_0,
	switches_in_export_1,
	switches_in_export_2,
	switches_in_export_3,
	switches_in_export_4,
	switches_in_export_5,
	switches_in_export_6,
	switches_in_export_7,
	switches_in_export_8,
	switches_in_export_9)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	readdata_0;
output 	readdata_1;
output 	readdata_2;
output 	readdata_3;
output 	readdata_4;
output 	readdata_5;
output 	readdata_6;
output 	readdata_7;
output 	readdata_8;
output 	readdata_9;
input 	int_nxt_addr_reg_dly_3;
input 	int_nxt_addr_reg_dly_2;
input 	clk_clk;
input 	switches_in_export_0;
input 	switches_in_export_1;
input 	switches_in_export_2;
input 	switches_in_export_3;
input 	switches_in_export_4;
input 	switches_in_export_5;
input 	switches_in_export_6;
input 	switches_in_export_7;
input 	switches_in_export_8;
input 	switches_in_export_9;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[1]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;
wire \read_mux_out[8]~combout ;
wire \read_mux_out[9]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\read_mux_out[8]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\read_mux_out[9]~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!switches_in_export_0),
	.datab(!int_nxt_addr_reg_dly_3),
	.datac(!int_nxt_addr_reg_dly_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h4040404040404040;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[1] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[7] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[8] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8] .extended_lut = "off";
defparam \read_mux_out[8] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[8] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[9] (
	.dataa(!int_nxt_addr_reg_dly_3),
	.datab(!int_nxt_addr_reg_dly_2),
	.datac(!switches_in_export_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[9] .extended_lut = "off";
defparam \read_mux_out[9] .lut_mask = 64'h0808080808080808;
defparam \read_mux_out[9] .shared_arith = "off";

endmodule
