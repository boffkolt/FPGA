
module niosii (
	buts_external_connection_export,
	clk_clk,
	leds_external_connection_export);	

	input	[7:0]	buts_external_connection_export;
	input		clk_clk;
	output	[7:0]	leds_external_connection_export;
endmodule
